module conv8_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [1024-1:0] input_act,
    output logic [1024-1:0] output_act,
    output logic ready
);

logic [1024-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 16'sd 20505) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6697) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27560) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4296) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13076) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10714) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26804) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11421) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28909) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3841) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19288) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23805) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14971) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7637) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19338) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30113) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10704) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11261) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15253) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8792) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22077) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29648) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2456) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24134) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21775) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9253) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20756) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28945) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6413) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29843) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28023) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18725) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13513) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4689) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29228) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7594) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31506) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19812) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23031) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3103) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18696) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9452) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12498) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4920) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32406) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22980) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10663) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1517) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10984) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18296) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27174) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25821) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17760) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19495) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20270) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18894) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9560) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16376) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12623) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7141) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6146) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21409) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24113) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_101[7:0]) +
	( 11'sd 686) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10761) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7638) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23969) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23038) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19888) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28606) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12254) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1765) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1119) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28755) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7476) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25875) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11241) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20187) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2485) * $signed(input_fmap_126[7:0]) +
	( 11'sd 973) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 13'sd 3136) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9039) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6374) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28531) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27408) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18260) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12164) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28290) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12683) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28834) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23510) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19719) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17815) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19616) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12895) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7230) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30166) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30090) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5054) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18206) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18330) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15879) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15687) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6323) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29761) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13815) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4665) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5133) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2859) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3992) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21543) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21694) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12181) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29997) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32596) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22190) * $signed(input_fmap_47[7:0]) +
	( 5'sd 14) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24693) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17217) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29495) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21054) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32632) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24330) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32437) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31968) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1452) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18560) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19525) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31062) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21652) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9291) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_69[7:0]) +
	( 11'sd 770) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2534) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28452) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31609) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7989) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_79[7:0]) +
	( 9'sd 207) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11656) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3868) * $signed(input_fmap_84[7:0]) +
	( 13'sd 4030) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8236) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27561) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9164) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10727) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31944) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8688) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15109) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25786) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17820) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9636) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31624) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7159) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28921) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9062) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24985) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22164) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25415) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22378) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19963) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27556) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13021) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_118[7:0]) +
	( 11'sd 643) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22103) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19653) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17551) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29269) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 16'sd 28115) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29871) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20896) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8401) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12574) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15373) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3787) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4426) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22642) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28279) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13720) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9516) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22243) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_14[7:0]) +
	( 5'sd 10) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22910) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19968) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28612) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30659) * $signed(input_fmap_19[7:0]) +
	( 11'sd 827) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17997) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26240) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26912) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15947) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3488) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28317) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11331) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13056) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1117) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9493) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_42[7:0]) +
	( 14'sd 8114) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16639) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_46[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8266) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16315) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10556) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13759) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18390) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18944) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23281) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30870) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7038) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30743) * $signed(input_fmap_62[7:0]) +
	( 10'sd 493) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30873) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20443) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32041) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31713) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7369) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16276) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29368) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6379) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31124) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21212) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8720) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2336) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20933) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21580) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13901) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13370) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5194) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_86[7:0]) +
	( 9'sd 164) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7792) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28118) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30450) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26440) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15349) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2846) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3096) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15779) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13364) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5045) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23082) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11670) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2065) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29362) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28974) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31666) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6347) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17959) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3640) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25402) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20769) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29302) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11444) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6312) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 16'sd 23679) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30705) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22098) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1243) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1075) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11580) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29494) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11104) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9247) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28754) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10371) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11132) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18158) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12267) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22903) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17899) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18713) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_26[7:0]) +
	( 10'sd 447) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14361) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29912) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21214) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21485) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20552) * $signed(input_fmap_33[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5087) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8923) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21041) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28894) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7753) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14206) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25549) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8880) * $signed(input_fmap_43[7:0]) +
	( 10'sd 376) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17557) * $signed(input_fmap_45[7:0]) +
	( 11'sd 614) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32511) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11768) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10731) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18280) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12670) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13395) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6992) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26012) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4100) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1640) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21371) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11371) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19881) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28259) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23376) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25545) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18841) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3202) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31622) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_71[7:0]) +
	( 11'sd 638) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24260) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25617) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3886) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27692) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14670) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26282) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2663) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1914) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22883) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18220) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17723) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24973) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13096) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21944) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17717) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13193) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28788) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1361) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3557) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25504) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18368) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20138) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10593) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4336) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5704) * $signed(input_fmap_107[7:0]) +
	( 11'sd 1002) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12737) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4413) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28716) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21504) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25551) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27625) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14777) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23320) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7538) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 16'sd 19104) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1607) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19756) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1246) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32539) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31783) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26033) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17494) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13847) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_11[7:0]) +
	( 14'sd 8161) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7648) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8741) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23956) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_21[7:0]) +
	( 11'sd 544) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20741) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26309) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_28[7:0]) +
	( 11'sd 894) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1790) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23215) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30427) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27826) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9640) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14160) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5718) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29441) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7460) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14979) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27987) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21077) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21028) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19881) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19192) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26205) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3372) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27689) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6473) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13650) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14035) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22521) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18979) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5643) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21290) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21371) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32450) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30076) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7732) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22395) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30850) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7560) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26428) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8802) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10044) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31663) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5264) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1255) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28211) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12816) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23238) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16763) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11884) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4668) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8560) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26502) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_100[7:0]) +
	( 10'sd 354) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4449) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32121) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25088) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19441) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10693) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24759) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7423) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5970) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2633) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13830) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29693) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29602) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16148) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6783) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8197) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11331) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_125[7:0]) +
	( 11'sd 783) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 14'sd 5222) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13043) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17091) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19691) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20607) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23493) * $signed(input_fmap_10[7:0]) +
	( 13'sd 4028) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13112) * $signed(input_fmap_12[7:0]) +
	( 11'sd 734) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10367) * $signed(input_fmap_14[7:0]) +
	( 11'sd 619) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1782) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8105) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10579) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11175) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24686) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21797) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26171) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32274) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17025) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13915) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4878) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27970) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8278) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14546) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25196) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9765) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22074) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17069) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11679) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27483) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4583) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2207) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13268) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28030) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8226) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2698) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8253) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29476) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9738) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12346) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18382) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7336) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26685) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25058) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6241) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2219) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25138) * $signed(input_fmap_83[7:0]) +
	( 10'sd 396) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14571) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3531) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13168) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6368) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8529) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3684) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18584) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6906) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25311) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5290) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24973) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19959) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10938) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26367) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2944) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19041) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16464) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10223) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31751) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17618) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23294) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15414) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26346) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29663) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12713) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8921) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14899) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 16'sd 22718) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12365) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_4[7:0]) +
	( 12'sd 2040) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25742) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15442) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7727) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14261) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24269) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27860) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12560) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18706) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19242) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31279) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26841) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29425) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16013) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3330) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9174) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20482) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26561) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29771) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19401) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32235) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25573) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13809) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22727) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7986) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30069) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3168) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15392) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17030) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25366) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7204) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23122) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28707) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29766) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25921) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9332) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13792) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11686) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8758) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28256) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18564) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10240) * $signed(input_fmap_69[7:0]) +
	( 11'sd 601) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26625) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30718) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31768) * $signed(input_fmap_76[7:0]) +
	( 11'sd 721) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13933) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9962) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21495) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14021) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16313) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26066) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4747) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19659) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1220) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4104) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7902) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11567) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20053) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10487) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31901) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17669) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23834) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13037) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3500) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21476) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29735) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26549) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21212) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23669) * $signed(input_fmap_112[7:0]) +
	( 11'sd 638) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28670) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26693) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3579) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10639) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11375) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29999) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_123[7:0]) +
	( 10'sd 284) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31503) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29164) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5021) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 14'sd 4468) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14848) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8267) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12167) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18588) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1032) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31515) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17924) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25850) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22318) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22151) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1693) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30775) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14833) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3579) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31982) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12519) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28348) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8492) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1678) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1453) * $signed(input_fmap_26[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19764) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15112) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26638) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26386) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5249) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18804) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26086) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9235) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7709) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11057) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31070) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24090) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32011) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17964) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26421) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32124) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19973) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12196) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20244) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17025) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28403) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24847) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14949) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22215) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24193) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13154) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9464) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17401) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27656) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22747) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5282) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16283) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18372) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11829) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3000) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7828) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27061) * $signed(input_fmap_95[7:0]) +
	( 10'sd 475) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6609) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9252) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26486) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30288) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27031) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8701) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11608) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18961) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22069) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10219) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22514) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8875) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5507) * $signed(input_fmap_117[7:0]) +
	( 9'sd 147) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21253) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1692) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32750) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23160) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12354) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22353) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7992) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 16'sd 23721) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14619) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16425) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4443) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17882) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10596) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14129) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14691) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22762) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21905) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28192) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31621) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21312) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16848) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22138) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25035) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24992) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14124) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1247) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8792) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18594) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5039) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29732) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22120) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23904) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20731) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20433) * $signed(input_fmap_34[7:0]) +
	( 10'sd 413) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7656) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12100) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26273) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4840) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20975) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6847) * $signed(input_fmap_42[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7733) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11135) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1441) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25667) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16096) * $signed(input_fmap_50[7:0]) +
	( 13'sd 4046) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15620) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24198) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15894) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19762) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16968) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24082) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15718) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26193) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21325) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13110) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17702) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15655) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17520) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30967) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16160) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18915) * $signed(input_fmap_85[7:0]) +
	( 13'sd 4014) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20256) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24538) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29720) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21665) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23297) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27257) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10444) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17595) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2821) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28092) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32091) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7421) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18993) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22728) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11090) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2543) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5197) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25258) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19547) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12336) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6532) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18775) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29752) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23535) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19509) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 16'sd 23827) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24258) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14082) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23065) * $signed(input_fmap_3[7:0]) +
	( 10'sd 461) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3359) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18044) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23390) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27112) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28851) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31855) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30306) * $signed(input_fmap_13[7:0]) +
	( 11'sd 634) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4115) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10530) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31894) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_20[7:0]) +
	( 10'sd 441) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26482) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20862) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18205) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20601) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25774) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6676) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22512) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27649) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4986) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24923) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20576) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4227) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22922) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8368) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13980) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19432) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12653) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13906) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20340) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27765) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28314) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21432) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23957) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16605) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11250) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9014) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11253) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9664) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29142) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5045) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5851) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21696) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21080) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2728) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9925) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14913) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22377) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21895) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20865) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30462) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5829) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18383) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1291) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1468) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27073) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16768) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29610) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4656) * $signed(input_fmap_94[7:0]) +
	( 7'sd 40) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31171) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13652) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1870) * $signed(input_fmap_99[7:0]) +
	( 11'sd 795) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28324) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5671) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1710) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30976) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20322) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25145) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11715) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21039) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29442) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17707) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14606) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8750) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9015) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13361) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9533) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26121) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28163) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9394) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1733) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23549) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 16'sd 20998) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1917) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4762) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20482) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20289) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14419) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27168) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8668) * $signed(input_fmap_9[7:0]) +
	( 11'sd 781) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31811) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27212) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15796) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24472) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5248) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20871) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12275) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19135) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18987) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2218) * $signed(input_fmap_27[7:0]) +
	( 11'sd 747) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30876) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15138) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5522) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18154) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9474) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7097) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17245) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5988) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20634) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31825) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15635) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21069) * $signed(input_fmap_47[7:0]) +
	( 10'sd 282) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30706) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6945) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4511) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19643) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15585) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23920) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7080) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15629) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_59[7:0]) +
	( 8'sd 109) * $signed(input_fmap_60[7:0]) +
	( 11'sd 633) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18071) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13940) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32184) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23694) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17802) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5273) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16477) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18962) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27695) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27822) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22296) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5144) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5354) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5550) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27444) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7296) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30603) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1982) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29418) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20567) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13972) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7992) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10007) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29251) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9180) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8558) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28691) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27767) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19837) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6207) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20101) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2093) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21369) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2425) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24818) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25641) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21660) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19869) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28766) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30057) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8582) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11694) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 16'sd 26626) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5690) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9587) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8717) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21854) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29493) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22570) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24423) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14979) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26677) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29142) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31348) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25913) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11571) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25742) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31798) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31018) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29731) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14180) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13610) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2377) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8654) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22551) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24050) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31790) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4341) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26254) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27540) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11589) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32064) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22565) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12512) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5207) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2594) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9727) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21551) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12267) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15545) * $signed(input_fmap_63[7:0]) +
	( 11'sd 517) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25753) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14177) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14665) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9746) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20302) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27222) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11143) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18576) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4937) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13046) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28747) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16414) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27674) * $signed(input_fmap_85[7:0]) +
	( 11'sd 989) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1536) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14555) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12068) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21736) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22460) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1904) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22418) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1852) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5792) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30476) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30358) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32031) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1114) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23279) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8066) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1749) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28736) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30253) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18824) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20658) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15845) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8077) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8960) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23748) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9782) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32754) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31683) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8425) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 16'sd 22130) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5826) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6761) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27017) * $signed(input_fmap_3[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12829) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_6[7:0]) +
	( 14'sd 8102) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2460) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19028) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5570) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29929) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27863) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20218) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16022) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7768) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15619) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27707) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9032) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16494) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30440) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30879) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23153) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16967) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2048) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27592) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23353) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6967) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7207) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19012) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30018) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19674) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10873) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2048) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2362) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8853) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26514) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3266) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11077) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1201) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27127) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30905) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29396) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30862) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9091) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26785) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11054) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15881) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27674) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8754) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23462) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7993) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12351) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2537) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23184) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16442) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12150) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28161) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25472) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6132) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11825) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15587) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31034) * $signed(input_fmap_94[7:0]) +
	( 12'sd 2025) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3554) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16099) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18664) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13279) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6778) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17239) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15412) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16956) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14100) * $signed(input_fmap_110[7:0]) +
	( 7'sd 39) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26406) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3440) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19128) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6784) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19799) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 12'sd 1615) * $signed(input_fmap_0[7:0]) +
	( 11'sd 558) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2833) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32085) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_9[7:0]) +
	( 11'sd 536) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16448) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20165) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23473) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28924) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17640) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19218) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25092) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5463) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14230) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12573) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6362) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9819) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20871) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30369) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25908) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21512) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2185) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11881) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29333) * $signed(input_fmap_40[7:0]) +
	( 11'sd 881) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24450) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26733) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19289) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14957) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24420) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24073) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15280) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32111) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21922) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25558) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14122) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24495) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14053) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10416) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15886) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30981) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30177) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13405) * $signed(input_fmap_68[7:0]) +
	( 15'sd 16371) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15928) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27986) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16074) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11313) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32684) * $signed(input_fmap_76[7:0]) +
	( 8'sd 85) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21479) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15032) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14750) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21003) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30987) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10917) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12735) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17804) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16835) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30967) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25915) * $signed(input_fmap_100[7:0]) +
	( 11'sd 660) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4479) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30611) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17227) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12157) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16329) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24272) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18113) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5043) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25587) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17428) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20055) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29925) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19336) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_121[7:0]) +
	( 12'sd 2001) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7316) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30695) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17533) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 15'sd 15306) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18608) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31648) * $signed(input_fmap_2[7:0]) +
	( 11'sd 620) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7481) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20268) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20980) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6735) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17085) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14558) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6231) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23038) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5881) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2869) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30235) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25033) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16180) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12808) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3109) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6524) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5809) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_31[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15348) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8700) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19346) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20431) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1771) * $signed(input_fmap_38[7:0]) +
	( 8'sd 65) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25193) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27921) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22872) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10455) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7414) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30605) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4210) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30348) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2390) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9851) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18088) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14992) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3061) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22610) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2180) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25526) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12644) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17260) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23114) * $signed(input_fmap_77[7:0]) +
	( 10'sd 466) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31650) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19997) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11981) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2887) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8638) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7056) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18358) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28225) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2724) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7477) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26011) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1850) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4445) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27967) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19328) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13826) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19381) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10534) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22847) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28731) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29566) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24004) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25420) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4683) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17580) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1858) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2406) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3605) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2432) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4477) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13219) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16183) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 14'sd 4429) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32758) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19998) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32522) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11754) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26253) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2509) * $signed(input_fmap_14[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28954) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13516) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18090) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22481) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14287) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31232) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19539) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22051) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5092) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1397) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26204) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26169) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12107) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20605) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14909) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6333) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2646) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6618) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9963) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29654) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31839) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16398) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13813) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10821) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13778) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26989) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21221) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7909) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20390) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27500) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5639) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21747) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5554) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1817) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4187) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14642) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6140) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6714) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14935) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25330) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31437) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20261) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10554) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6987) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28039) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8266) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23908) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21688) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3674) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26605) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29319) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4475) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25120) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28349) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9348) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11656) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5826) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10130) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21392) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6674) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21325) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14305) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27192) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28690) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2614) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10885) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19031) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22689) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10657) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30507) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15265) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 16'sd 21863) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22443) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10363) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18441) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17633) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22461) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5442) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8634) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28499) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13521) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8775) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12821) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18656) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11222) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25785) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1579) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2524) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25797) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8718) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19089) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26591) * $signed(input_fmap_24[7:0]) +
	( 11'sd 695) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4728) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21536) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4304) * $signed(input_fmap_31[7:0]) +
	( 9'sd 156) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23380) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24358) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7374) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2621) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15515) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4857) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20528) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5260) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23671) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5109) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30860) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15628) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22523) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7240) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29443) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27676) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27662) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20420) * $signed(input_fmap_62[7:0]) +
	( 10'sd 478) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12004) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29236) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23129) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16771) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16661) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10727) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4623) * $signed(input_fmap_77[7:0]) +
	( 10'sd 303) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5076) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12849) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16171) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22744) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30841) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_91[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23285) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3654) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31891) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6910) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22176) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29874) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13479) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10867) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32738) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23871) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23411) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22710) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17104) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5276) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13371) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8163) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28685) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7899) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16377) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9486) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9907) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11465) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16158) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 16'sd 20135) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3252) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13784) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24786) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16543) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32626) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20898) * $signed(input_fmap_10[7:0]) +
	( 10'sd 298) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3122) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17537) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22853) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32113) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26748) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15622) * $signed(input_fmap_20[7:0]) +
	( 11'sd 568) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9315) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29579) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8365) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29537) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14291) * $signed(input_fmap_28[7:0]) +
	( 11'sd 931) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12207) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7286) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17785) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28986) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15347) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32517) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10532) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8563) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_40[7:0]) +
	( 10'sd 434) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24518) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22930) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20137) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31604) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17465) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6395) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24131) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23262) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11471) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6201) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7810) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20501) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20129) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30977) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9248) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18562) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26699) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22224) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27594) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15459) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2775) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24995) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9766) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7187) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4212) * $signed(input_fmap_87[7:0]) +
	( 11'sd 827) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18886) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28896) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2631) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28621) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13518) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2989) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1293) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10821) * $signed(input_fmap_97[7:0]) +
	( 11'sd 578) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6431) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30062) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21428) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30797) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8341) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17164) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29590) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17879) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4971) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28198) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6271) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16090) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 15'sd 8495) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4411) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18664) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27865) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22676) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19125) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2411) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31566) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4734) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13138) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29218) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14067) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25351) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10828) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31191) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_28[7:0]) +
	( 11'sd 887) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12209) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25484) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4149) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9157) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29006) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10998) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3655) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31629) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17035) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30062) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10753) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5692) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9420) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4382) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22297) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28090) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25138) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20578) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16745) * $signed(input_fmap_54[7:0]) +
	( 11'sd 526) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11912) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30004) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1552) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21041) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16861) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10602) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8820) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5408) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24448) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3518) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13680) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30059) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20820) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14911) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16290) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8701) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31752) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10397) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15870) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14462) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25652) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2493) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31233) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18030) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31431) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8439) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15054) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8847) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17615) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15576) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4520) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2588) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5341) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7668) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22997) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22046) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2170) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14949) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7339) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17865) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22051) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26751) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31566) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32106) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13449) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28287) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32037) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11799) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29200) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 15'sd 8365) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23428) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18475) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32192) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1944) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19100) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13056) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17330) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3427) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13737) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18274) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17694) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25522) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17186) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26692) * $signed(input_fmap_23[7:0]) +
	( 11'sd 851) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22493) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7830) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15467) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27798) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17236) * $signed(input_fmap_33[7:0]) +
	( 11'sd 512) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24808) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29703) * $signed(input_fmap_37[7:0]) +
	( 11'sd 760) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17881) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26723) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15054) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18291) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3829) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6952) * $signed(input_fmap_45[7:0]) +
	( 11'sd 856) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27220) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14275) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6355) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16401) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2202) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13510) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21696) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28435) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23106) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3573) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10271) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4317) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10521) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29916) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23875) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28568) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29645) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2123) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4615) * $signed(input_fmap_79[7:0]) +
	( 11'sd 832) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17490) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6039) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3623) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18801) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24737) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19641) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9385) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31559) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5218) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2495) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27762) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20581) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13818) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21583) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8778) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15967) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4104) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30541) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22575) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17335) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13797) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16509) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3855) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28576) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4790) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32098) * $signed(input_fmap_123[7:0]) +
	( 8'sd 90) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30180) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 16'sd 30915) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29520) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15340) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19205) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21400) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19070) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15677) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5305) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17969) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23507) * $signed(input_fmap_10[7:0]) +
	( 14'sd 8127) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17216) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8866) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30833) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22162) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8576) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25603) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26972) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32430) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14341) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14241) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26197) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27028) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31348) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29303) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25339) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7785) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17973) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30344) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9087) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26864) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17421) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21164) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22396) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26635) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6182) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2787) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14748) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25824) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13847) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20819) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3258) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17321) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17641) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6038) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10884) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13737) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14884) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26379) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4423) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19912) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3875) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17920) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11363) * $signed(input_fmap_75[7:0]) +
	( 9'sd 188) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29959) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10499) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24370) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20725) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21049) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4764) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9479) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7554) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2771) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9876) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11107) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19302) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_96[7:0]) +
	( 11'sd 1013) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5138) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16119) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29624) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24949) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5005) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7947) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9087) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8935) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24432) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18417) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6863) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31153) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23135) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4849) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23073) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5181) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5887) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29569) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32760) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4343) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11373) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 13'sd 3306) * $signed(input_fmap_0[7:0]) +
	( 11'sd 907) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32646) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10327) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28784) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29372) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8123) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20806) * $signed(input_fmap_9[7:0]) +
	( 7'sd 49) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14907) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27245) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15895) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18745) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29135) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6473) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32520) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1225) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24861) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19858) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29337) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27141) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15612) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30047) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11800) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29902) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16949) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13682) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10358) * $signed(input_fmap_34[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28173) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22716) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27200) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25258) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29119) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26804) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4258) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32628) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15418) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21426) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20665) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9661) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5757) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17606) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10169) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30600) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7089) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6222) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13646) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22011) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12688) * $signed(input_fmap_67[7:0]) +
	( 14'sd 8101) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3105) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1125) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14234) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10594) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9310) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23447) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_79[7:0]) +
	( 10'sd 430) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3165) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9804) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20442) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17750) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1085) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25021) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11336) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29437) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8248) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7984) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15225) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10346) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11257) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19471) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7417) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18763) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25966) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20839) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11243) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15762) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25819) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11577) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19619) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5322) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9524) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26078) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8819) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5495) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 14'sd 5402) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14022) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25016) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30291) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27411) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14205) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11892) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2269) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29218) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19629) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27935) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13909) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24543) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29945) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20267) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23706) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17263) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30588) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28791) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3943) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11228) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15610) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6657) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8351) * $signed(input_fmap_30[7:0]) +
	( 10'sd 280) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5311) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11018) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6441) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2077) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18198) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30548) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5908) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8481) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27402) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4546) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2340) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11705) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26518) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28158) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30847) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2096) * $signed(input_fmap_54[7:0]) +
	( 10'sd 308) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19817) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14873) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19286) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8237) * $signed(input_fmap_60[7:0]) +
	( 11'sd 982) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_63[7:0]) +
	( 11'sd 804) * $signed(input_fmap_64[7:0]) +
	( 7'sd 33) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22861) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21598) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17562) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12941) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14757) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32552) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27913) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10218) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14651) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17415) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13509) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21145) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2353) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2667) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27287) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5807) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25833) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14604) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24394) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15084) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3572) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26004) * $signed(input_fmap_101[7:0]) +
	( 10'sd 447) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8605) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12839) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20234) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1377) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9588) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19942) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_112[7:0]) +
	( 11'sd 652) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14718) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10299) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7066) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4626) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7740) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20709) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27199) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 13'sd 4055) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2588) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12084) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26723) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19088) * $signed(input_fmap_5[7:0]) +
	( 10'sd 436) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21895) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26265) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5584) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14569) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18805) * $signed(input_fmap_13[7:0]) +
	( 11'sd 901) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7505) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17908) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5309) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15222) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14210) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16167) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18592) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13838) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9510) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27332) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1042) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3122) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2259) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19454) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5307) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24519) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10979) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23109) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9412) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15900) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23825) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12850) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19660) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_52[7:0]) +
	( 11'sd 614) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20402) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32584) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19992) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_59[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6514) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32388) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13104) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31897) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3041) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19244) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26036) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8488) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21436) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30433) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31053) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5895) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25519) * $signed(input_fmap_83[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17756) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26835) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4371) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7270) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2482) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8729) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14995) * $signed(input_fmap_92[7:0]) +
	( 4'sd 5) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28948) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20567) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14030) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9447) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28419) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22832) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12984) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3859) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12266) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_107[7:0]) +
	( 11'sd 915) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21174) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17743) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3073) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22813) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18509) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12388) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15445) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11065) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25276) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19276) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6597) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25972) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25945) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_124[7:0]) +
	( 11'sd 628) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10703) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18577) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 14'sd 4331) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26021) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26466) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23467) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8097) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11593) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31574) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28274) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28395) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8504) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23853) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19971) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23073) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30833) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32346) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10692) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24343) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18724) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27829) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15424) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30942) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19521) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25242) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22070) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3813) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9981) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3747) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1081) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24110) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_48[7:0]) +
	( 11'sd 911) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14777) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8483) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23157) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28644) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23944) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7105) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_60[7:0]) +
	( 12'sd 2031) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27160) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6079) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11936) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6585) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1224) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19348) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21319) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6042) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2637) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23802) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6948) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19755) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2508) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30468) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9851) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25415) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8412) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5054) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20753) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27383) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24752) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1410) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23814) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9891) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26366) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8981) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17237) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17373) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29721) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27155) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25667) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25925) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11577) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10553) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27713) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8002) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2928) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9437) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6884) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16445) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7222) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13628) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 16'sd 21030) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27701) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18418) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19509) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28049) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28684) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13315) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14903) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29476) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11164) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14742) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23948) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21479) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24887) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6557) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4610) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7207) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28817) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11706) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15436) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5261) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28993) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30065) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20556) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20653) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20844) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24909) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29375) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_39[7:0]) +
	( 6'sd 27) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6687) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15248) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3138) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11888) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18609) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18522) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23279) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12394) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22855) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19716) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28458) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18244) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4987) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23225) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16254) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21236) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_64[7:0]) +
	( 11'sd 544) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15683) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21393) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24599) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29147) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29836) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18677) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3475) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19764) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8789) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19982) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30136) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28611) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31498) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3699) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5503) * $signed(input_fmap_88[7:0]) +
	( 9'sd 199) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14177) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29536) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25147) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18468) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28944) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30468) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13696) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19021) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7641) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17624) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5794) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19094) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_104[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22502) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5415) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31209) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26489) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26297) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10337) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10189) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7985) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31821) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27383) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20905) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8958) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 14'sd 7289) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28540) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30851) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1154) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22252) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8792) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_7[7:0]) +
	( 9'sd 135) * $signed(input_fmap_8[7:0]) +
	( 8'sd 84) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22106) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31231) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22066) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18197) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24859) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8707) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20066) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18399) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19958) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22215) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20703) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20159) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13410) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17065) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14127) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4845) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14359) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29945) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23633) * $signed(input_fmap_39[7:0]) +
	( 10'sd 291) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27806) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32408) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2503) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1610) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27512) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1335) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30217) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26973) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9960) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20404) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18205) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12629) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18822) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20185) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4171) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10050) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3620) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5942) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1938) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27108) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21216) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27275) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16938) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20969) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13092) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12063) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25160) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18809) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16649) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22355) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27842) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18615) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2321) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19205) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23185) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1225) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2861) * $signed(input_fmap_96[7:0]) +
	( 9'sd 227) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31852) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21856) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4519) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5273) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26295) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14789) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17793) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16363) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6809) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25688) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1942) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10707) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5179) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29028) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15681) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28630) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5516) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27101) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5284) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20482) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 16'sd 16825) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6589) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28252) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17158) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23209) * $signed(input_fmap_6[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10059) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30510) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12397) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19765) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30002) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30363) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_18[7:0]) +
	( 10'sd 487) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5476) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32677) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7869) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8280) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20242) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20757) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25323) * $signed(input_fmap_35[7:0]) +
	( 11'sd 959) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2123) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4666) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30276) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28567) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15634) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4916) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14680) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23074) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26906) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2757) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29114) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15723) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21487) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17260) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16980) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26796) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9833) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28046) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12741) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18342) * $signed(input_fmap_69[7:0]) +
	( 11'sd 819) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15572) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29411) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28075) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29292) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14275) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25491) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9861) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5325) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15533) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3052) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25421) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25286) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16877) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18574) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14447) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10149) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15254) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6105) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3394) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25442) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25492) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29182) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19725) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23358) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30833) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6855) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16230) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12546) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31909) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20343) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2317) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31998) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22038) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30225) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16143) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21910) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11453) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27292) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17843) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 16'sd 32254) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10265) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5994) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16467) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29960) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5246) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7187) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20715) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30417) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1290) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31233) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3869) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15163) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2833) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13919) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22392) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_20[7:0]) +
	( 11'sd 771) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8123) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15245) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7838) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29515) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23084) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9325) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9786) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10716) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29985) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14383) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25826) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9104) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9427) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25822) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28522) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27967) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22606) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11297) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12958) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24982) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24156) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13837) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29735) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18712) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6247) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3253) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6534) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20712) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23947) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14808) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9450) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4970) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13548) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5720) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10215) * $signed(input_fmap_77[7:0]) +
	( 10'sd 258) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31236) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23038) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24315) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20156) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26039) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26090) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1307) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28896) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27731) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28505) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16690) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14412) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12147) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7845) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8724) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15167) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16027) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16313) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_109[7:0]) +
	( 11'sd 654) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6164) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22741) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9171) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_115[7:0]) +
	( 11'sd 746) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2418) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14949) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11333) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19135) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32393) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4807) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10123) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31679) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24039) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 16'sd 30888) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22061) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10068) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10982) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16718) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_7[7:0]) +
	( 11'sd 756) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29051) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1863) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9676) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24567) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4182) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7925) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23332) * $signed(input_fmap_21[7:0]) +
	( 11'sd 650) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32353) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27737) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3731) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8349) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9243) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14970) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24767) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26485) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4948) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6735) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24229) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7198) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29532) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10297) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11766) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29248) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12595) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_54[7:0]) +
	( 5'sd 14) * $signed(input_fmap_55[7:0]) +
	( 10'sd 322) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14067) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17264) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_61[7:0]) +
	( 11'sd 562) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6091) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31787) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2195) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21817) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25616) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32564) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27806) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17016) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1366) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8023) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12190) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7097) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23616) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31087) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23900) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10409) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21728) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25554) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16889) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24308) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12009) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18551) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28077) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5601) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14031) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9234) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17290) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31765) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1426) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14867) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16097) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26525) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23713) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11408) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29669) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31771) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24098) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17373) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7016) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4560) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27274) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24268) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23626) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22226) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32664) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27251) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22531) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26812) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21035) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 16'sd 25727) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17498) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15669) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12401) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18309) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10482) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2806) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9010) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27161) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28019) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1853) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30659) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11517) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27435) * $signed(input_fmap_21[7:0]) +
	( 11'sd 582) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20115) * $signed(input_fmap_23[7:0]) +
	( 11'sd 933) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18940) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11013) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4696) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5259) * $signed(input_fmap_29[7:0]) +
	( 11'sd 930) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7054) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15363) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11872) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20037) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19549) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29240) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13012) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27039) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30231) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26803) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13771) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22045) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29117) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29092) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18929) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13300) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24585) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26049) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26838) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30747) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19436) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4409) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14614) * $signed(input_fmap_65[7:0]) +
	( 11'sd 732) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25914) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30863) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15598) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8431) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22070) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12567) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8222) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27738) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4148) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29919) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16324) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19490) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9181) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27244) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20533) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1992) * $signed(input_fmap_92[7:0]) +
	( 10'sd 288) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19264) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14293) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32627) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26107) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4675) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28787) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28144) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29118) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27767) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8875) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7085) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16560) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25536) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15785) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9521) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20495) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24928) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27369) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21026) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19651) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18254) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3831) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 15'sd 9549) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18046) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4238) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24423) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15349) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12649) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18922) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7906) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24236) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_11[7:0]) +
	( 11'sd 884) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4626) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6523) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31616) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21721) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24993) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24627) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18373) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31439) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10962) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14710) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14082) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21252) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23167) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8334) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22722) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5670) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30822) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14378) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30434) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27743) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16969) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13558) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12087) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7170) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18372) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28993) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27188) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31328) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28883) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29412) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23164) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24953) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27474) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31367) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24198) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6164) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13950) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5588) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6166) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32432) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17883) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27365) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9663) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14988) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6081) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3731) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5810) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7430) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6843) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29068) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25590) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2855) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14555) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8695) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2813) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19850) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13620) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22061) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32617) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18523) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1061) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22970) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29121) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31742) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20546) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12237) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14227) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14585) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32394) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 15'sd 9763) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24897) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19706) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20431) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1422) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22989) * $signed(input_fmap_6[7:0]) +
	( 11'sd 626) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21949) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4126) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17522) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7011) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23758) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12466) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3837) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21295) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6348) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14450) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26612) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24714) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21968) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4834) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28342) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7364) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22106) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5619) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29384) * $signed(input_fmap_32[7:0]) +
	( 8'sd 78) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17760) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31827) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27222) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3965) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20023) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14185) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1082) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11183) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9763) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6886) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8495) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1936) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19623) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20025) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19074) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28366) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26647) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15103) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18865) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5741) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25871) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14433) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16673) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9516) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22730) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10539) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10170) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30274) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3658) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25910) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13655) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19279) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9687) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6352) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28115) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3494) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31819) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15212) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32570) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28336) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30460) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12248) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12629) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1267) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24903) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7326) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15219) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11945) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17933) * $signed(input_fmap_114[7:0]) +
	( 9'sd 252) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18225) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6884) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5226) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11585) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 16'sd 21689) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13051) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21595) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16981) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28678) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20704) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31515) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18445) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28952) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16701) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7972) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28837) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_18[7:0]) +
	( 11'sd 606) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29109) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_21[7:0]) +
	( 10'sd 504) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8803) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5665) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19415) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32088) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5098) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30265) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23885) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12906) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17868) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28446) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13797) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3331) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29777) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27162) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4872) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20639) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20799) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29231) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11597) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6456) * $signed(input_fmap_57[7:0]) +
	( 14'sd 8031) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26584) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9560) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23546) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5617) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9123) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4839) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32012) * $signed(input_fmap_68[7:0]) +
	( 15'sd 16119) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12501) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12733) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24234) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15052) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11401) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22415) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12175) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20389) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1137) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2939) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26970) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3231) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30641) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27101) * $signed(input_fmap_95[7:0]) +
	( 11'sd 577) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8751) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27983) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13960) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5651) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10246) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7396) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5465) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3385) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16431) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5411) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4797) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9842) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18594) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18892) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8378) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10778) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16922) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3813) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14639) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6341) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 16'sd 21931) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9402) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10748) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26414) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5050) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4202) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16281) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12556) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29821) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3179) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25738) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30895) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1456) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9498) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12934) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28493) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21557) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26484) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27171) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18519) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16045) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17641) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9813) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1591) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23850) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18337) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21594) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18541) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31507) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4211) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22277) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8017) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1292) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18424) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22059) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17394) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9888) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22597) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30591) * $signed(input_fmap_54[7:0]) +
	( 9'sd 252) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7645) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6266) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15868) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21113) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9626) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13457) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24644) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9488) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20039) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21368) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32184) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29164) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20518) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14411) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13998) * $signed(input_fmap_81[7:0]) +
	( 9'sd 198) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29251) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15967) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29706) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9651) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13838) * $signed(input_fmap_95[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29765) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31867) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20251) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28361) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17046) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10282) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12334) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17824) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16424) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20481) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22271) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8992) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31814) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30231) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1551) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5776) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6551) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21428) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26820) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_122[7:0]) +
	( 10'sd 327) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16090) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 14'sd 7179) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26451) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9691) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12772) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29096) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2103) * $signed(input_fmap_7[7:0]) +
	( 8'sd 91) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21687) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29837) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9114) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29462) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6999) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11303) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30638) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4341) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26251) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18475) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12872) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9961) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4622) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7982) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30613) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16887) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9877) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17058) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29713) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15709) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23285) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15461) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20038) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17866) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26477) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6076) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15415) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13243) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1042) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10712) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7830) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11201) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30881) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11881) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16587) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9456) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22134) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27603) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12809) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21794) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27946) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16279) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22821) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23172) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10829) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21720) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18088) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5353) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13206) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13858) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23836) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7752) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15429) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27922) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22279) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21880) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18629) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1903) * $signed(input_fmap_101[7:0]) +
	( 11'sd 694) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18204) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21874) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20499) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7372) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26942) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10876) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32156) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20282) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32653) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16944) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5951) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4713) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24256) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27224) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3139) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22497) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19597) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6857) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5284) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1769) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 14'sd 7507) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12435) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20015) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25129) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18376) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16220) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1098) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9821) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3903) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14980) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1842) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25246) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9467) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23195) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21877) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29528) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27052) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22450) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26906) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23087) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21126) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23294) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23124) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7478) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7891) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29451) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21268) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29252) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10205) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16604) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2351) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16461) * $signed(input_fmap_52[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19064) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23063) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27365) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27731) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5692) * $signed(input_fmap_63[7:0]) +
	( 11'sd 602) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16855) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9956) * $signed(input_fmap_67[7:0]) +
	( 11'sd 762) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15144) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20588) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27696) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23432) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5182) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15631) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20289) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15740) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22888) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28069) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8484) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31766) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27339) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5674) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26023) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7368) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23878) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_93[7:0]) +
	( 11'sd 730) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14639) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25615) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29632) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7126) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12498) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10009) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20130) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22422) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5492) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1221) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28855) * $signed(input_fmap_116[7:0]) +
	( 11'sd 643) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13468) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11306) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30289) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3347) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6460) * $signed(input_fmap_126[7:0]) +
	( 10'sd 302) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 16'sd 30216) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6799) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29557) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21397) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2266) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20759) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29212) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7479) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13395) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31840) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31576) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3757) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31592) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25045) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5934) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10370) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1328) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24140) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19110) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19924) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24514) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30559) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6140) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12565) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25785) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7218) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17926) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11960) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16125) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16059) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31782) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9430) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29892) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16695) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12882) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9537) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19416) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32031) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7140) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28369) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26160) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1777) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32184) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6133) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24083) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28125) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26311) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5294) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2487) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10669) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10084) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5561) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30134) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27727) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22336) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2427) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23736) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19198) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15349) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21107) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4905) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15179) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26578) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13890) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21679) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16204) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18765) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6915) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3559) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29773) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10336) * $signed(input_fmap_111[7:0]) +
	( 11'sd 680) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12607) * $signed(input_fmap_113[7:0]) +
	( 14'sd 8015) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4945) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9805) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3578) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15868) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32165) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6286) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19379) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8236) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32026) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 16'sd 22755) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30597) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21270) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25298) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21680) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19230) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17891) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4493) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21650) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21290) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16404) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18291) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31493) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30927) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29650) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29644) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2289) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24208) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24122) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32100) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28345) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19022) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6270) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17801) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17507) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20814) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21100) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13165) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22853) * $signed(input_fmap_45[7:0]) +
	( 10'sd 272) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21448) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12300) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1236) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32243) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17989) * $signed(input_fmap_52[7:0]) +
	( 11'sd 933) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26091) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16822) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31930) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13046) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12063) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32028) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14502) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26586) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19530) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16637) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3355) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2563) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2855) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27759) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25679) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17067) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8379) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30560) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12921) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24440) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12904) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21061) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19488) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10824) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14728) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6219) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4347) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23439) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7505) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14474) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16842) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22463) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21763) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21035) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9068) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17589) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29417) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19852) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14289) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1896) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32292) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17299) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10270) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4506) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30848) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_121[7:0]) +
	( 11'sd 818) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7618) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24099) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10837) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 15'sd 9132) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15173) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14911) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13301) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18733) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25834) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3994) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28747) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26512) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17649) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23329) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10031) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14748) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9188) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4218) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8938) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8981) * $signed(input_fmap_23[7:0]) +
	( 14'sd 8009) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1410) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21804) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31805) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7975) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25585) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23118) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_35[7:0]) +
	( 9'sd 194) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19159) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25181) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5720) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13481) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7768) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4929) * $signed(input_fmap_42[7:0]) +
	( 10'sd 356) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2441) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20025) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6311) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14411) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18062) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26410) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10473) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8285) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28608) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19934) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10774) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18496) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18096) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5909) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12731) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3438) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3486) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13511) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26663) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17594) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24834) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12635) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4573) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13948) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18412) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3834) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15195) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17269) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31557) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23894) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11096) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22135) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22422) * $signed(input_fmap_94[7:0]) +
	( 10'sd 287) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4788) * $signed(input_fmap_96[7:0]) +
	( 11'sd 864) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25391) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18104) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32487) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29414) * $signed(input_fmap_106[7:0]) +
	( 11'sd 931) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24962) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22862) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16681) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3992) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27205) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_114[7:0]) +
	( 9'sd 178) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30488) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3367) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15889) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29346) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25779) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5828) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29513) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 13'sd 3646) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18181) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1908) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8684) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_5[7:0]) +
	( 11'sd 810) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30445) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12787) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6551) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19777) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_15[7:0]) +
	( 11'sd 813) * $signed(input_fmap_16[7:0]) +
	( 12'sd 2036) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22614) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3250) * $signed(input_fmap_24[7:0]) +
	( 7'sd 42) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29446) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8178) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28059) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20696) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25700) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23179) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24796) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16513) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10641) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6950) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7689) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21975) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11823) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27023) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24381) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1423) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29237) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4308) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23667) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22123) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26971) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28628) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8446) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22677) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11600) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10904) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6514) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8486) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6807) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4398) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19956) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6014) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4313) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30515) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13814) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10142) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17832) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18727) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24768) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32543) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14052) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3491) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3650) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26616) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14458) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15075) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29638) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17045) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15653) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11404) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8716) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5535) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29582) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10142) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10364) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5405) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15872) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_120[7:0]) +
	( 11'sd 771) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1995) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16384) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22146) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 14'sd 5210) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31753) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_5[7:0]) +
	( 11'sd 1018) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23062) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3974) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8560) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11333) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17511) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26934) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11137) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7405) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5903) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3397) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21624) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26464) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20551) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12418) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15256) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31382) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14758) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14963) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_38[7:0]) +
	( 11'sd 711) * $signed(input_fmap_39[7:0]) +
	( 11'sd 818) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29326) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18005) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12550) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7267) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6313) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9063) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_53[7:0]) +
	( 11'sd 616) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14084) * $signed(input_fmap_57[7:0]) +
	( 11'sd 759) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12442) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3269) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20578) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22136) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28622) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2687) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6521) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_66[7:0]) +
	( 11'sd 802) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_68[7:0]) +
	( 10'sd 279) * $signed(input_fmap_69[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7727) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29661) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20004) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19056) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18861) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21861) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12929) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10031) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2544) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4220) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25147) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9943) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13894) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15858) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9109) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17809) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2981) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13048) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29555) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17783) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3695) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17831) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14919) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10264) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21658) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31428) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21398) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6713) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5198) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10651) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7945) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27074) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5528) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16230) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_124[7:0]) +
	( 10'sd 431) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2502) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 16'sd 22319) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6030) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20009) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7565) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18740) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2094) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6567) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19836) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11470) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24761) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24083) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31201) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27337) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25876) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26450) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25597) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20542) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18577) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3789) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21528) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23809) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7467) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9381) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11100) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25675) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30622) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20356) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10071) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19792) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5651) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28522) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9050) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29422) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8695) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7130) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18387) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11728) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8006) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21990) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7747) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26502) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9428) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16370) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7529) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13488) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18010) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23427) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17700) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31544) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16812) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25800) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18148) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25244) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20571) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19610) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1858) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20181) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16283) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14038) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19903) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26128) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7170) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3169) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12114) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10891) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31854) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9881) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25218) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29304) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20640) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1426) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32724) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7477) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20388) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24979) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24293) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13046) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7645) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11781) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22043) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21782) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15610) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14903) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17302) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25219) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 16'sd 24719) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23860) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29793) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3165) * $signed(input_fmap_3[7:0]) +
	( 10'sd 305) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22977) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10214) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14470) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23088) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1913) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31524) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22254) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9411) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15076) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5324) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7162) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18874) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26840) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11080) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25488) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11912) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12613) * $signed(input_fmap_32[7:0]) +
	( 10'sd 304) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31369) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27653) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7490) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22947) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14083) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6574) * $signed(input_fmap_39[7:0]) +
	( 9'sd 221) * $signed(input_fmap_40[7:0]) +
	( 11'sd 855) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32712) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8623) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3945) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19151) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28907) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29415) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21210) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11952) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18397) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16098) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10663) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17303) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6799) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5320) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24759) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1399) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5874) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9688) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6594) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4553) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_68[7:0]) +
	( 10'sd 392) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11698) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6978) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24827) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6103) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6229) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1846) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16965) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20495) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30412) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19450) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23605) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26445) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4737) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15216) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6412) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26071) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19106) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22908) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4751) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8882) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9148) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6602) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20342) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10942) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20222) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18763) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4314) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32328) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3840) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18711) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20887) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29800) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27984) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3265) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20766) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 13'sd 2313) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29630) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9821) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_6[7:0]) +
	( 14'sd 8152) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9754) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29369) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27146) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3164) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22770) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19471) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30478) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11752) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21271) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8461) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2989) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_27[7:0]) +
	( 10'sd 353) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15367) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2861) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21712) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21538) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11376) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28116) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23352) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13870) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17228) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9492) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27152) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6786) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1230) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30126) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23636) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12706) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18930) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31627) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16140) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7970) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12108) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13328) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7856) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2685) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29443) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5088) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1216) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8829) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5835) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30422) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24144) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14670) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28403) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19978) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6496) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22309) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24630) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5504) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9317) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9791) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15249) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28296) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17376) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30437) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5744) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12234) * $signed(input_fmap_93[7:0]) +
	( 11'sd 686) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10449) * $signed(input_fmap_95[7:0]) +
	( 14'sd 8100) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5874) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19716) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4206) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17720) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4786) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9403) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15052) * $signed(input_fmap_105[7:0]) +
	( 11'sd 857) * $signed(input_fmap_106[7:0]) +
	( 14'sd 8011) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28958) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31943) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31986) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3112) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9709) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7333) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13041) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23733) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15906) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22443) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18274) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 16'sd 23370) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29715) * $signed(input_fmap_1[7:0]) +
	( 11'sd 883) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6597) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16677) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30985) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27323) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26203) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_14[7:0]) +
	( 9'sd 197) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10496) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4427) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21006) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15161) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25894) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6970) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9230) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29208) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17375) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31964) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3840) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28132) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25476) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15699) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19814) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_44[7:0]) +
	( 11'sd 554) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20613) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29657) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17156) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14234) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23326) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17866) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7034) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25248) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11432) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4272) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19027) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26557) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22666) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3104) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21176) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12871) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15278) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10767) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22698) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12064) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11060) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1727) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22413) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21415) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21134) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31305) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23615) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12522) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32720) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32094) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28945) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12777) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21341) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15816) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32719) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29154) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31826) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17065) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29553) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19327) * $signed(input_fmap_101[7:0]) +
	( 10'sd 409) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17795) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21612) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27090) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14202) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8896) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11945) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3171) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29665) * $signed(input_fmap_121[7:0]) +
	( 11'sd 890) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11546) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13378) * $signed(input_fmap_124[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22618) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 16'sd 25798) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19406) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1726) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22130) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7766) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30544) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6619) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15170) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8585) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13003) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3069) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27728) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7414) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26717) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28180) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18255) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20718) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11632) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17869) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6919) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6640) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3052) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16080) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16581) * $signed(input_fmap_41[7:0]) +
	( 9'sd 253) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21487) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26595) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5803) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29300) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13273) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3621) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7847) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6470) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7400) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3063) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31207) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9099) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31329) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6885) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13844) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17440) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22878) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1223) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14737) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10529) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1537) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20628) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1042) * $signed(input_fmap_76[7:0]) +
	( 10'sd 268) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12049) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31425) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15449) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26281) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_87[7:0]) +
	( 9'sd 150) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18280) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_90[7:0]) +
	( 11'sd 993) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23861) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27825) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6662) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5315) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3839) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2495) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28162) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7654) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23657) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27426) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31545) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12656) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2183) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3309) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23824) * $signed(input_fmap_114[7:0]) +
	( 12'sd 2031) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15264) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7310) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22353) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4889) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29284) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9463) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5585) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25116) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8657) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13913) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6108) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 16'sd 26259) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17258) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30276) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23769) * $signed(input_fmap_6[7:0]) +
	( 9'sd 213) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28011) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16208) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2848) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6739) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11653) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22232) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2887) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24525) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27660) * $signed(input_fmap_23[7:0]) +
	( 11'sd 695) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3969) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9934) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32674) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25115) * $signed(input_fmap_29[7:0]) +
	( 14'sd 8114) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12035) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22278) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31086) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5910) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6160) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24083) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17308) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12534) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5109) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_45[7:0]) +
	( 11'sd 885) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18318) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21599) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15648) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27153) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1207) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22729) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7241) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28806) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15129) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1889) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5704) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13382) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4375) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26163) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6111) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24160) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1636) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24534) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6466) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9077) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22068) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16807) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29457) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15699) * $signed(input_fmap_77[7:0]) +
	( 11'sd 592) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2050) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22172) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20532) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1463) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28780) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32712) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23511) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30369) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3315) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13500) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23897) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28415) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_99[7:0]) +
	( 11'sd 615) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32443) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11805) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31392) * $signed(input_fmap_105[7:0]) +
	( 11'sd 855) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16924) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8494) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15975) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19487) * $signed(input_fmap_112[7:0]) +
	( 11'sd 813) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32352) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13296) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13534) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14444) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25251) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 15'sd 13505) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26134) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12966) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26541) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14085) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30897) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11397) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_8[7:0]) +
	( 11'sd 736) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30391) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18382) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20533) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14808) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22752) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22251) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21389) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11736) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1572) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19391) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1154) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19921) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10391) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4446) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10362) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12002) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32711) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6105) * $signed(input_fmap_39[7:0]) +
	( 9'sd 133) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32692) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22022) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8804) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12564) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27750) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20277) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10082) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13972) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6071) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3036) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13940) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3182) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1048) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8627) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1243) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12380) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18290) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29363) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24398) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25334) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29354) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1696) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21232) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22167) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18145) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3603) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20388) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29562) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11656) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19360) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18829) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1074) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27395) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2237) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3013) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19063) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9608) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2922) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20376) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_114[7:0]) +
	( 11'sd 660) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26914) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21999) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17633) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21078) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14082) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4311) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18749) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 16'sd 29393) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10881) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32522) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5159) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32022) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7411) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30238) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29885) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21391) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22650) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15935) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32460) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22723) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9491) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28721) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1453) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26907) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26572) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20777) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21133) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15814) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5728) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28399) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11001) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27212) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14456) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13593) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13229) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22607) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21221) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20528) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8871) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8997) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6079) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29057) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31876) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15427) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32074) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19260) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12639) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19372) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2467) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17435) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13283) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22150) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6375) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5800) * $signed(input_fmap_69[7:0]) +
	( 10'sd 465) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25223) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12510) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6194) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21886) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7908) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31674) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22037) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28871) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8488) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22492) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11951) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26440) * $signed(input_fmap_88[7:0]) +
	( 13'sd 4030) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14149) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19506) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4433) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7730) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21061) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12035) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13602) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13053) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27039) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27910) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26026) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28263) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5497) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2482) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29369) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15283) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10415) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11377) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30730) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30038) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27361) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31386) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18208) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1129) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8825) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 14'sd 6203) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24841) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15655) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9215) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31650) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9237) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24600) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19933) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17878) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32236) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5612) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20889) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26149) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26788) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17267) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21009) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27590) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30764) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19019) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30094) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21658) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20364) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13110) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12523) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8710) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29374) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14006) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30888) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29470) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11400) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26822) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19869) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28491) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17400) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7784) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30699) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22817) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11206) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28628) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31979) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29093) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17062) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25462) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13146) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31273) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31955) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13378) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19717) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25415) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8777) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31097) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26045) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7141) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9798) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16112) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26729) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12340) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7532) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24778) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14692) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7203) * $signed(input_fmap_93[7:0]) +
	( 11'sd 969) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10061) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29306) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14404) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31194) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12379) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27804) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27524) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10755) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_108[7:0]) +
	( 11'sd 787) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5365) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2071) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24354) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14427) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32595) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26119) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13495) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_123[7:0]) +
	( 11'sd 982) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11349) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7192) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3630) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 16'sd 32187) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15195) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3935) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24505) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18270) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20948) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1554) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30695) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28856) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14180) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12043) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10884) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6837) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7272) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3090) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32431) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23410) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31145) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10533) * $signed(input_fmap_29[7:0]) +
	( 14'sd 8168) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10161) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6518) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21996) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4369) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28597) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27726) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11815) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9478) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7323) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3426) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27147) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18774) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2791) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18860) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10433) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_52[7:0]) +
	( 10'sd 386) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14179) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26564) * $signed(input_fmap_58[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20272) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12138) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16973) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25595) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22300) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4511) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18652) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23049) * $signed(input_fmap_76[7:0]) +
	( 8'sd 100) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21361) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10415) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18958) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29327) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32584) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11020) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5036) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1259) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29226) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6123) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2653) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10492) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32670) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29211) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19500) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7618) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7374) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22286) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15039) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10362) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3291) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2359) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17603) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15109) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9782) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13956) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16439) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19682) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10138) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8806) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19147) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24995) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14543) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10987) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 16'sd 26296) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14262) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15329) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4437) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9246) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12384) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1929) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8479) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12329) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5616) * $signed(input_fmap_20[7:0]) +
	( 11'sd 726) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10662) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12756) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2373) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30599) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29956) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16604) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28649) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17855) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31838) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21008) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29925) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12241) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12722) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22157) * $signed(input_fmap_45[7:0]) +
	( 11'sd 594) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32632) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1705) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21740) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19976) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6274) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4481) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30595) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26258) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31597) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26353) * $signed(input_fmap_60[7:0]) +
	( 9'sd 157) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25782) * $signed(input_fmap_62[7:0]) +
	( 9'sd 173) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14141) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3924) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24640) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24430) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11758) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25844) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25284) * $signed(input_fmap_71[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12832) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28222) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9696) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19155) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9450) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25396) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18201) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22555) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11397) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25459) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21751) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25004) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14830) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7086) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15283) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4855) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3651) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14224) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1549) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8340) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17628) * $signed(input_fmap_107[7:0]) +
	( 11'sd 689) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25551) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6390) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18907) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13520) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19685) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4637) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30419) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27865) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28760) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1431) * $signed(input_fmap_125[7:0]) +
	( 10'sd 461) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23173) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 16'sd 17852) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1534) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21869) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17853) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1700) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20818) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_8[7:0]) +
	( 11'sd 525) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18197) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19812) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7308) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31956) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_17[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1659) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4752) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31037) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31528) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1257) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28051) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14868) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19521) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2130) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17559) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4094) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16875) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30652) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17698) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11231) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13564) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8192) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23783) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2139) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28563) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18721) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21650) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31588) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15508) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28936) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7521) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1930) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25679) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22370) * $signed(input_fmap_60[7:0]) +
	( 11'sd 926) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23910) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23646) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20910) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24554) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25160) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28723) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6194) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18660) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23494) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3474) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25948) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28632) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14624) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14812) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6059) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27727) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8658) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17908) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22696) * $signed(input_fmap_87[7:0]) +
	( 11'sd 754) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15759) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18518) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5105) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10921) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13870) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20309) * $signed(input_fmap_97[7:0]) +
	( 11'sd 584) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19198) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31377) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_102[7:0]) +
	( 11'sd 708) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_104[7:0]) +
	( 13'sd 4056) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12244) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21278) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18938) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14362) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23483) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13783) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1827) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4318) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22096) * $signed(input_fmap_121[7:0]) +
	( 11'sd 785) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14018) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29580) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11009) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26785) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 16'sd 26575) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4114) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17090) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21298) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30128) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15233) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31959) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32312) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1861) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12090) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19674) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24341) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14672) * $signed(input_fmap_13[7:0]) +
	( 11'sd 725) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3646) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12486) * $signed(input_fmap_16[7:0]) +
	( 10'sd 275) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20921) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21456) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23566) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10902) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17593) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14337) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19910) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20472) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30536) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8591) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10925) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7144) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18223) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8661) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25281) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1467) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7439) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4599) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25114) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19385) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31973) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7860) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20368) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23410) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17557) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28460) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23067) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16015) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25593) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15764) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16805) * $signed(input_fmap_64[7:0]) +
	( 11'sd 660) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2147) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11455) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23733) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10422) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25285) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8643) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20298) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11608) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27386) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32527) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22741) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28266) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32375) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7652) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30968) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22767) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3142) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31627) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1876) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16142) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31278) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15996) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11473) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16200) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4321) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9516) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25920) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30498) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_117[7:0]) +
	( 12'sd 2032) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25915) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6897) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25753) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8386) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4839) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1858) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 15'sd 8304) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1622) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2358) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16329) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9555) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10705) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17091) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32098) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27094) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23196) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_11[7:0]) +
	( 9'sd 255) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2406) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20355) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27909) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23260) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4498) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16070) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22488) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6449) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20420) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6908) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20154) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13991) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30004) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20630) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8878) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18147) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31794) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18647) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13614) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16792) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12715) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17616) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24753) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2165) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23513) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21474) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31781) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32069) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15901) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30104) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2810) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3784) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23713) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23215) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30582) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22097) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12129) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4937) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1474) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_80[7:0]) +
	( 9'sd 209) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7582) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29700) * $signed(input_fmap_85[7:0]) +
	( 10'sd 383) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32049) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5425) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3593) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13737) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21871) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24939) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27006) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30025) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10523) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9235) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11879) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5112) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1900) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8385) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18284) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26712) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14730) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21419) * $signed(input_fmap_118[7:0]) +
	( 9'sd 138) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24918) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21237) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_122[7:0]) +
	( 11'sd 935) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24378) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30348) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11357) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 15'sd 11458) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7567) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27561) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12896) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10044) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12722) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30004) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18258) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12501) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12753) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29620) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26609) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19217) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19492) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2899) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21509) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4502) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27671) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1122) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15236) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6939) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21139) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24913) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19346) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17031) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6471) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20475) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31731) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6448) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30092) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28520) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3477) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32467) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1293) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22416) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11057) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22264) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25208) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13906) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14061) * $signed(input_fmap_63[7:0]) +
	( 10'sd 301) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26612) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21501) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21687) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22770) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13267) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31850) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30008) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18987) * $signed(input_fmap_76[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10550) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6278) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29501) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14927) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13472) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30523) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25631) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16816) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5695) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9147) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16748) * $signed(input_fmap_99[7:0]) +
	( 10'sd 491) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27817) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23032) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31990) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4583) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11110) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29414) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31694) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27913) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24643) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28490) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7695) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11809) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11949) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30561) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21890) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21711) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10977) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 16'sd 26653) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27728) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5825) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31831) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28785) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2093) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17445) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8494) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25369) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30105) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14004) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25121) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_22[7:0]) +
	( 11'sd 802) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4929) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5429) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16308) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31787) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3660) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3632) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30941) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32152) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10889) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14766) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22681) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31265) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28949) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18580) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3734) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14443) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23995) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26884) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21782) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23560) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25064) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15838) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12652) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10415) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11735) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12033) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28679) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26341) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5018) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22912) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28596) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29491) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31792) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30904) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_83[7:0]) +
	( 10'sd 300) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_85[7:0]) +
	( 11'sd 1020) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28723) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13565) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11473) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20193) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15348) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14796) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29664) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13709) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8935) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23313) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5636) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7361) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15374) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30754) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24208) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17532) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5163) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22562) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7329) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23793) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6568) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27081) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 14'sd 6025) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19535) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24363) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8017) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2798) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31159) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10761) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8513) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27455) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4572) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3897) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6333) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25622) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14634) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29507) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24716) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22584) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4862) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18121) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_31[7:0]) +
	( 13'sd 4060) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29464) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12660) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10756) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6884) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12865) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28504) * $signed(input_fmap_39[7:0]) +
	( 9'sd 225) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29922) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8004) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24738) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1675) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28792) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_51[7:0]) +
	( 9'sd 229) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5210) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25607) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3862) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28185) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12573) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26976) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15588) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15843) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11846) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10661) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11046) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11268) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14843) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10104) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28982) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2200) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23843) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10690) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12650) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25254) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7296) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27464) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15139) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17775) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17604) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9576) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13122) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_99[7:0]) +
	( 9'sd 150) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32209) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6670) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9471) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30502) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15021) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2303) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26550) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30181) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7597) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16969) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6430) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27315) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1302) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 16'sd 26662) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13195) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1976) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8729) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8218) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15060) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25968) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5514) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21035) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22438) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23360) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6349) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8429) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26189) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22408) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26134) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17824) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28289) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23293) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6401) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1029) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10928) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31164) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14150) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14648) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9154) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19158) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30873) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30469) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8552) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6615) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5527) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25303) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24460) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11379) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1656) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15472) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14322) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_55[7:0]) +
	( 11'sd 954) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24856) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22802) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5132) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31535) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9025) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14278) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13749) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16021) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5478) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20824) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24150) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25347) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9366) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28076) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31460) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22842) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24401) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26919) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29464) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20706) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2143) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31312) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4406) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1066) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15823) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26622) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_89[7:0]) +
	( 11'sd 724) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26214) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25307) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16434) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3788) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24631) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12730) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21815) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14329) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10741) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19951) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_104[7:0]) +
	( 11'sd 836) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29518) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10303) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1945) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1676) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9121) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5678) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31790) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29895) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29725) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23481) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8729) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25525) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6240) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 15'sd 8567) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8994) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4814) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6108) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10987) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10955) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9663) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17432) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24460) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16987) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28138) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21476) * $signed(input_fmap_19[7:0]) +
	( 8'sd 107) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23097) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9315) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16362) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7389) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6958) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8964) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11750) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14019) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13915) * $signed(input_fmap_37[7:0]) +
	( 10'sd 338) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15279) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28857) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23466) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32034) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9953) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28773) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6807) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9006) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17614) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31822) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14092) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15699) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3272) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31253) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8862) * $signed(input_fmap_57[7:0]) +
	( 13'sd 4084) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24781) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1983) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11156) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24406) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10594) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23540) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16287) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21358) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18161) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30748) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11750) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9130) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17361) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13895) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30080) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12048) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32179) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30957) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3731) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22098) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1875) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8460) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24937) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9655) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5001) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19500) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28097) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24582) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14854) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28708) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1329) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15054) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7902) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28774) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12074) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13643) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6362) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26785) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4893) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2306) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10307) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1193) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20138) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 15'sd 15178) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14338) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3510) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20984) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12040) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10401) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9235) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11412) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16816) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3239) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12475) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28359) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6001) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8399) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17087) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_18[7:0]) +
	( 11'sd 761) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23439) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31200) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27048) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4828) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7206) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28183) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13187) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5731) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1657) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26556) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21267) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16240) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24711) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9661) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20582) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30195) * $signed(input_fmap_44[7:0]) +
	( 9'sd 226) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2957) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14949) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23597) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3994) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21054) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11130) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9978) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4621) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17150) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20458) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19875) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16059) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20305) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12917) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1916) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6632) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25131) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26280) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11037) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27010) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2540) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3695) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6134) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10598) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28490) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27445) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3085) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5855) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1168) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30056) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10518) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2318) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28182) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18844) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12225) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14115) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2906) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11237) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15565) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22244) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18922) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3494) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31721) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2759) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11371) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26693) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10156) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7982) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6510) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25882) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6956) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4834) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18462) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29348) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 15'sd 14178) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31813) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1555) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24836) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11297) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21131) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31489) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31974) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17700) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12114) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25662) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23278) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32473) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20553) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8469) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15680) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13609) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32546) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7765) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_29[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13597) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10596) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12535) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11489) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17392) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23620) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14093) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6821) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1137) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11864) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21215) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25283) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29499) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13724) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6596) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7339) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27481) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1343) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32491) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10679) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7470) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13012) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28848) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14030) * $signed(input_fmap_69[7:0]) +
	( 11'sd 766) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26246) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21902) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_77[7:0]) +
	( 11'sd 849) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_79[7:0]) +
	( 11'sd 949) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_81[7:0]) +
	( 7'sd 58) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25177) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7968) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7576) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12830) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6880) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32362) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17386) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10136) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_100[7:0]) +
	( 7'sd 38) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28260) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22448) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2777) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1633) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3146) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26700) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2299) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26288) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12569) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8710) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25093) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21944) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17716) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19196) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28949) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3691) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2682) * $signed(input_fmap_124[7:0]) +
	( 8'sd 109) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11658) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20183) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 15'sd 9899) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28787) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29081) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23285) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19709) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2402) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12745) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8016) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18759) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27181) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28244) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18910) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30756) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21539) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25463) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6866) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16878) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23139) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6427) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3504) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4649) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29534) * $signed(input_fmap_38[7:0]) +
	( 10'sd 298) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25269) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12151) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27817) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25613) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31303) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11234) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22397) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29269) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5598) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8019) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12452) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31903) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13721) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29729) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24676) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8675) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31102) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10498) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13459) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30061) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3448) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22826) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31751) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6978) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32306) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14302) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22825) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19369) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14257) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5910) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9108) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21788) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8751) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14172) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2817) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15753) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9329) * $signed(input_fmap_103[7:0]) +
	( 12'sd 2021) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32059) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6009) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32230) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28502) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19843) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5711) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3785) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28482) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28529) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7856) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14281) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27314) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 16'sd 21566) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11539) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5528) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1250) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_6[7:0]) +
	( 11'sd 537) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29783) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1119) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4706) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14599) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18584) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23760) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10192) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19510) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11011) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28146) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5983) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3055) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18277) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23125) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2904) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2501) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17622) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27344) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22831) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17384) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5221) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30436) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14553) * $signed(input_fmap_39[7:0]) +
	( 6'sd 20) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25593) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1871) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14818) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7009) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17869) * $signed(input_fmap_49[7:0]) +
	( 13'sd 4083) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1988) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29200) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8738) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11876) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6910) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8415) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23535) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17903) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3640) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25177) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18129) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32343) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5348) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27750) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12236) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6762) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16673) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29217) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16917) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11801) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18932) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24430) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1287) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16832) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2089) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31646) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29646) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14655) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26052) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_99[7:0]) +
	( 9'sd 238) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5486) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30116) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21185) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22932) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21347) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4694) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25675) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27762) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26112) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15997) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10498) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20893) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24617) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7218) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31309) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21805) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 16'sd 16551) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7540) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26016) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7187) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22941) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8497) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31976) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15868) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16565) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13859) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27794) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29504) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13537) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3030) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26754) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4207) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21839) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10463) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13273) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17205) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11619) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11492) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25678) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_44[7:0]) +
	( 10'sd 282) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30896) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2573) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26578) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7501) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4169) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3030) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6016) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26189) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24378) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_60[7:0]) +
	( 9'sd 180) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25907) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20549) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18451) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15635) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2646) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22009) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25739) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10865) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15296) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16971) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29092) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9963) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21146) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14831) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_86[7:0]) +
	( 10'sd 425) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4483) * $signed(input_fmap_88[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10546) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11109) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25281) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4132) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28779) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3666) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24104) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22963) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19229) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26279) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24391) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11176) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30232) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22579) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9612) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30282) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30808) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1925) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13405) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29780) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16861) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12506) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15190) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28158) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13848) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12366) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27230) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 13'sd 3799) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25301) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13924) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26079) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9918) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_7[7:0]) +
	( 11'sd 806) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20311) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11147) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16772) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23653) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26285) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2278) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6233) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14118) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29942) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23747) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22357) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11886) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12239) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5020) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7513) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10100) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20846) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21723) * $signed(input_fmap_33[7:0]) +
	( 11'sd 793) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15893) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21009) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13950) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4884) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19264) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15263) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25131) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19579) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2810) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20605) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6448) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20670) * $signed(input_fmap_50[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10389) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1657) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11679) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16652) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22448) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29305) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29574) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15303) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22736) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17085) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17586) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17298) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31994) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18820) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13755) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13617) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17901) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21195) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9359) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15130) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28339) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31100) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3881) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17075) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6429) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31861) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3826) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9216) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12309) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30342) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25199) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5662) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21618) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20008) * $signed(input_fmap_108[7:0]) +
	( 11'sd 901) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7437) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28802) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13191) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5028) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5247) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17664) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21478) * $signed(input_fmap_122[7:0]) +
	( 11'sd 521) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17182) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14711) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31312) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16347) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 14'sd 5892) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18545) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21564) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19603) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5105) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7775) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6268) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25702) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_12[7:0]) +
	( 11'sd 930) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16588) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29501) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7278) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20926) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24910) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12688) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16692) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16922) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3932) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12229) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27007) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10031) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26855) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21546) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26740) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28903) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4552) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19733) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10967) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13889) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22171) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16835) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16853) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15533) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2921) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23755) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8199) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30357) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_58[7:0]) +
	( 10'sd 266) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7051) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6631) * $signed(input_fmap_61[7:0]) +
	( 11'sd 683) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16442) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3334) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19123) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10287) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31368) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14989) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24863) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27558) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15893) * $signed(input_fmap_73[7:0]) +
	( 9'sd 145) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3622) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13237) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4776) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22780) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7343) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32137) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5289) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1063) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3781) * $signed(input_fmap_89[7:0]) +
	( 12'sd 2000) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3128) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8395) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26309) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26242) * $signed(input_fmap_96[7:0]) +
	( 11'sd 668) * $signed(input_fmap_97[7:0]) +
	( 10'sd 435) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32059) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31912) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11408) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32180) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10573) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14052) * $signed(input_fmap_108[7:0]) +
	( 10'sd 354) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30391) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14572) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25062) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7616) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3627) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9159) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8887) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14183) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9414) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2922) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31728) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30232) * $signed(input_fmap_125[7:0]) +
	( 10'sd 442) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23583) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 15'sd 11500) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12253) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7657) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23834) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25543) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23281) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17961) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11694) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27586) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21421) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12594) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11653) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3800) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9642) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27977) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19465) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11553) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27719) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3040) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17330) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1777) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2199) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27245) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24577) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25736) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28722) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30701) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12364) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16725) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29966) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14797) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24472) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2968) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23215) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18655) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6770) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28846) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19771) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25672) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1149) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3634) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13705) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13049) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29124) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18563) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9307) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7220) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32539) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12495) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7771) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21743) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7916) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21243) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_80[7:0]) +
	( 11'sd 569) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12181) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_84[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15931) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13481) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10904) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25995) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24262) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12614) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17994) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18302) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4400) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28471) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12680) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16138) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8971) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3442) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28875) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29902) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27680) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4256) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12468) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5702) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4488) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1348) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2687) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 16'sd 25132) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6428) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10522) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7360) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_6[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21152) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18288) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22175) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13996) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16374) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22080) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27749) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23983) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2729) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25896) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29971) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3443) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26088) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6253) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_34[7:0]) +
	( 14'sd 8111) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2468) * $signed(input_fmap_38[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31792) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4246) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23372) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10734) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24141) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9924) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7506) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4951) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13819) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10111) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17794) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16695) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10991) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26116) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31976) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4246) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30097) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18457) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30830) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21805) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7849) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_73[7:0]) +
	( 11'sd 952) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8210) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13077) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28458) * $signed(input_fmap_80[7:0]) +
	( 10'sd 280) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21090) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22764) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13809) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17565) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16725) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25388) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6515) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19337) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27857) * $signed(input_fmap_96[7:0]) +
	( 10'sd 429) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11210) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12676) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8669) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15032) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25846) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17468) * $signed(input_fmap_104[7:0]) +
	( 11'sd 535) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23611) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19290) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11472) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27354) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20396) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21528) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12185) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7747) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12896) * $signed(input_fmap_119[7:0]) +
	( 11'sd 964) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2240) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17465) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21099) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12948) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6124) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1981) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 16'sd 20716) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13160) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22811) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25416) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19306) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26050) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19843) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21948) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29329) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22169) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27716) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32726) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12172) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3583) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4217) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10887) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17286) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16402) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1185) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1636) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27127) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18136) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29884) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20718) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4175) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6182) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4187) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13939) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28513) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3588) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23835) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6925) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15292) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19768) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29953) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2609) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32088) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_60[7:0]) +
	( 9'sd 219) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15587) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27724) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14337) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9840) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4136) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31092) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13547) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12927) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27152) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18165) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6061) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25081) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16029) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3637) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18927) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10203) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8500) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20507) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22865) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9166) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_91[7:0]) +
	( 10'sd 510) * $signed(input_fmap_92[7:0]) +
	( 11'sd 930) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29116) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30455) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32298) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20301) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11748) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30083) * $signed(input_fmap_101[7:0]) +
	( 8'sd 64) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_106[7:0]) +
	( 14'sd 8063) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1556) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22824) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23319) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30650) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25121) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19819) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7874) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12394) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21952) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25566) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1794) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18308) * $signed(input_fmap_124[7:0]) +
	( 13'sd 4040) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26019) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 16'sd 17200) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25900) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17731) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6739) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25814) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32368) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24353) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18933) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22407) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21739) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27084) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6823) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19010) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11703) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21358) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27346) * $signed(input_fmap_16[7:0]) +
	( 11'sd 752) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6225) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23858) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21282) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4603) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1363) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14927) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16449) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3154) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2083) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21329) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18958) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25589) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27368) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8376) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1572) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31711) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7533) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24517) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20194) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3142) * $signed(input_fmap_48[7:0]) +
	( 11'sd 856) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30498) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9247) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32588) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31589) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15445) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31715) * $signed(input_fmap_56[7:0]) +
	( 11'sd 766) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18636) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8980) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19713) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23759) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7446) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13726) * $signed(input_fmap_67[7:0]) +
	( 14'sd 8017) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1535) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30797) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8757) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27023) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17759) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15391) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4468) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18348) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10540) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15424) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16031) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11070) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21175) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7158) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4933) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4543) * $signed(input_fmap_91[7:0]) +
	( 11'sd 793) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24002) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24956) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14946) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21524) * $signed(input_fmap_100[7:0]) +
	( 11'sd 891) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12623) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11310) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12240) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17502) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32689) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30273) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25591) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_115[7:0]) +
	( 10'sd 430) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4783) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22653) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9812) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8187) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18922) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24004) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14213) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22071) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 15'sd 11691) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28347) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30793) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11007) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5349) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12953) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27109) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5757) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15311) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1894) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6761) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12483) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4890) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19100) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13287) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31740) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24827) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24104) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6936) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22877) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22204) * $signed(input_fmap_31[7:0]) +
	( 11'sd 881) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19914) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9355) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31946) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1125) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31599) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26302) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31441) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26364) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7206) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24783) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22811) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11912) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32358) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25040) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29128) * $signed(input_fmap_55[7:0]) +
	( 9'sd 217) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29582) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10126) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27414) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_62[7:0]) +
	( 11'sd 993) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24431) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8571) * $signed(input_fmap_65[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10928) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5294) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6195) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31599) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15427) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4987) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5966) * $signed(input_fmap_73[7:0]) +
	( 13'sd 4008) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30187) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2679) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10737) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9664) * $signed(input_fmap_78[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28348) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15111) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2779) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13832) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21902) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23916) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6836) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20767) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29372) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5785) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30116) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27613) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2829) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6274) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_96[7:0]) +
	( 3'sd 3) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27470) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18530) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2185) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6950) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27345) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28846) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24996) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31078) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13483) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26709) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16637) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21982) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7720) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6466) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13969) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18918) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7038) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28952) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27485) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 16'sd 31952) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29017) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6879) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_3[7:0]) +
	( 11'sd 577) * $signed(input_fmap_4[7:0]) +
	( 9'sd 170) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3256) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29274) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4365) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27872) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28286) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24605) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_15[7:0]) +
	( 10'sd 379) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8802) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4558) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3334) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23571) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10127) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28674) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28058) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17236) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19241) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30416) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16357) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32052) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30514) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8281) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28047) * $signed(input_fmap_39[7:0]) +
	( 13'sd 4083) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26866) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18169) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18186) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13423) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19546) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26408) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27668) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31028) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5559) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14744) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1828) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12248) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19822) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19546) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15390) * $signed(input_fmap_62[7:0]) +
	( 10'sd 291) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4611) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9114) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22542) * $signed(input_fmap_66[7:0]) +
	( 12'sd 2012) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7041) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9044) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14333) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27918) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15539) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16263) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6114) * $signed(input_fmap_81[7:0]) +
	( 11'sd 793) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3713) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25921) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10915) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5390) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5910) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11968) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21448) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15778) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24265) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10789) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8799) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30723) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1176) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7444) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1574) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5419) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21669) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15993) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3059) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29159) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28085) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16662) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27259) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7509) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15050) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5761) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11669) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27174) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30037) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21064) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28761) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 16'sd 24246) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10773) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7924) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28499) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5427) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26013) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14911) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26340) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23088) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32000) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7158) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15118) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31112) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18669) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2670) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26668) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22091) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16499) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24359) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25374) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17120) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22118) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27751) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10487) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1915) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6068) * $signed(input_fmap_45[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9434) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18780) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12664) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29557) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24696) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25669) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24682) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22524) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21159) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13193) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17038) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17320) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11693) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20929) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3414) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16324) * $signed(input_fmap_75[7:0]) +
	( 11'sd 1002) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9427) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1064) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31777) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32481) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2814) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8164) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13417) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12071) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10607) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23125) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12483) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3314) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13827) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24790) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18747) * $signed(input_fmap_103[7:0]) +
	( 10'sd 346) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18663) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24745) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5332) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29320) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29821) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11918) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25401) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18955) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10806) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11084) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10654) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32095) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14253) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21154) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15664) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8597) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20564) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7882) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 16'sd 17614) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24783) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29610) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14502) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24859) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8095) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2303) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11355) * $signed(input_fmap_11[7:0]) +
	( 8'sd 79) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2114) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32170) * $signed(input_fmap_14[7:0]) +
	( 10'sd 422) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22698) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1961) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1745) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5179) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15516) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30614) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27704) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30146) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10894) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5517) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26733) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18260) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4947) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29383) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1616) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12522) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10156) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32573) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31146) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20595) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4474) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30323) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24405) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6733) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25814) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23367) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4591) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22847) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27073) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_61[7:0]) +
	( 10'sd 340) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4880) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7621) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6996) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31389) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32338) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3315) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1278) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21322) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4538) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19463) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32235) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8498) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29005) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23252) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23224) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10068) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26570) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1197) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22643) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29261) * $signed(input_fmap_95[7:0]) +
	( 11'sd 535) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26790) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8334) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30863) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15266) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6551) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5268) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31037) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14430) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8647) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25769) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19812) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6929) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7577) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23371) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15402) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22994) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17970) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27807) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24600) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 15'sd 9322) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22657) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21821) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21517) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32512) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8654) * $signed(input_fmap_8[7:0]) +
	( 11'sd 662) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4373) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32694) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25296) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5303) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14134) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23820) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10927) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4308) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1911) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27181) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5761) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28511) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21638) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27524) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28243) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18474) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7593) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12110) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26747) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1731) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15748) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6665) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9078) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7195) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4381) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9943) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12232) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16064) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13830) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29258) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13785) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6372) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_63[7:0]) +
	( 11'sd 672) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4379) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16383) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21362) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19844) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3590) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27601) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23473) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11414) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8530) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6357) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6279) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23334) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30587) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15764) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_85[7:0]) +
	( 11'sd 532) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1118) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20615) * $signed(input_fmap_90[7:0]) +
	( 11'sd 887) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12567) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9198) * $signed(input_fmap_93[7:0]) +
	( 11'sd 690) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23293) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29532) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23575) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22044) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10706) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8633) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14556) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28253) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24752) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16016) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5750) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20678) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1228) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30749) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5431) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7942) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25565) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5107) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22760) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 15'sd 12584) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28322) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31023) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18542) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23735) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17640) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16721) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30191) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19150) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6069) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24461) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31022) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6896) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29646) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5917) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6911) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13746) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9234) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15039) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13360) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13335) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32488) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13312) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27992) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16752) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28274) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27845) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16586) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11449) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22958) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28241) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29379) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23587) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29328) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14768) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16089) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13934) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21633) * $signed(input_fmap_58[7:0]) +
	( 10'sd 325) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20757) * $signed(input_fmap_60[7:0]) +
	( 10'sd 490) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19814) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25064) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29285) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17831) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14484) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14010) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29764) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21642) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30393) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30138) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13829) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20006) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_82[7:0]) +
	( 11'sd 583) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26047) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21347) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29449) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21462) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23675) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31399) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15302) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24497) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2938) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20042) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26465) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12153) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2248) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14163) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17653) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7451) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28052) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6012) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4834) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6714) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14059) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19965) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19908) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18618) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27183) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6528) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30831) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 15'sd 12441) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10191) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2492) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25795) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23393) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11293) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19868) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8875) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21191) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3390) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23263) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24037) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6629) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10737) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18409) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21900) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22241) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3879) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14375) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22621) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9497) * $signed(input_fmap_25[7:0]) +
	( 9'sd 182) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5324) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25714) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21237) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11091) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22143) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25935) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10290) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31490) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5243) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22668) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30686) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5834) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28496) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18148) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32409) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32041) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19727) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5754) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10908) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28565) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28173) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21518) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31994) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22066) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13783) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10093) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22095) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5085) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11408) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10385) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17157) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6980) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30569) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25268) * $signed(input_fmap_80[7:0]) +
	( 11'sd 935) * $signed(input_fmap_81[7:0]) +
	( 9'sd 133) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24688) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11609) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30042) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31854) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5047) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6465) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1224) * $signed(input_fmap_96[7:0]) +
	( 11'sd 991) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1549) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15132) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4549) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1336) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3349) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16435) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11240) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14687) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23835) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25983) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10423) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2388) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26213) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22472) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_123[7:0]) +
	( 10'sd 338) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 15'sd 15539) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22813) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29146) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9829) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27766) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4723) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14002) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19257) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25932) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14982) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23961) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28612) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20347) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11631) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23033) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23335) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27343) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25127) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28440) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19013) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31674) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14873) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23597) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6079) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16197) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16002) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26947) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9542) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8330) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28802) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31586) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29766) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24722) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15879) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31571) * $signed(input_fmap_55[7:0]) +
	( 11'sd 835) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22511) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8691) * $signed(input_fmap_58[7:0]) +
	( 10'sd 442) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15188) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28362) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6679) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5736) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12027) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27405) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17276) * $signed(input_fmap_69[7:0]) +
	( 11'sd 915) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21504) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20158) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10025) * $signed(input_fmap_73[7:0]) +
	( 11'sd 567) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32204) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15478) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19208) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25113) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9574) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8938) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19756) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19991) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11493) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32718) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15572) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27083) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4935) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20810) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24661) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22983) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24759) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_99[7:0]) +
	( 10'sd 357) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9578) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22332) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14114) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28792) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25881) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1084) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27350) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15427) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11380) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13095) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24770) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6852) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32363) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12552) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 15'sd 15648) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2745) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29460) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17297) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_7[7:0]) +
	( 8'sd 65) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6886) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13568) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28367) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19073) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18625) * $signed(input_fmap_15[7:0]) +
	( 11'sd 514) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21140) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7681) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17963) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8678) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30701) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9548) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31421) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25904) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22234) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29852) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24535) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25993) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17928) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3680) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27524) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29912) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20566) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3723) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22671) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9706) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20987) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_56[7:0]) +
	( 12'sd 2044) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13657) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18759) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7922) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21917) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30692) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7229) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29982) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25657) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13248) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28804) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20330) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32073) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13423) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1062) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18696) * $signed(input_fmap_83[7:0]) +
	( 11'sd 649) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24220) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8765) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26379) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14094) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23931) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13149) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31162) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31133) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17464) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27455) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21114) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5597) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23209) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29969) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20474) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30204) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3771) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14878) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8750) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15068) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22980) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23353) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11129) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6718) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9709) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22159) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4595) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 15'sd 12365) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22257) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20433) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1984) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8258) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22955) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1981) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5837) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7095) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32392) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19621) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23248) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11586) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32730) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19727) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23034) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21627) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22272) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11148) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4340) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25645) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23856) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26910) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4044) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22710) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2947) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5698) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17572) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15852) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3364) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3418) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12991) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21780) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10957) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17204) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5418) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28328) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23783) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7500) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9070) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27894) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16065) * $signed(input_fmap_58[7:0]) +
	( 10'sd 266) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11441) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6669) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_62[7:0]) +
	( 9'sd 187) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17049) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22276) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5367) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22322) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26424) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27282) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16203) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10003) * $signed(input_fmap_73[7:0]) +
	( 13'sd 4094) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4495) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2311) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30526) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26479) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2364) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26546) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15293) * $signed(input_fmap_83[7:0]) +
	( 10'sd 341) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17966) * $signed(input_fmap_85[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28578) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22852) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32430) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1372) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16190) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21041) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28884) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19970) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16774) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9879) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3762) * $signed(input_fmap_101[7:0]) +
	( 10'sd 309) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23043) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24405) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18987) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25589) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10477) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12340) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22116) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23938) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3982) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13688) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18405) * $signed(input_fmap_118[7:0]) +
	( 10'sd 311) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27759) * $signed(input_fmap_120[7:0]) +
	( 11'sd 765) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19021) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29973) * $signed(input_fmap_125[7:0]) +
	( 10'sd 295) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20383) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 11'sd 527) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31071) * $signed(input_fmap_1[7:0]) +
	( 11'sd 606) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23826) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6538) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29732) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25684) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25569) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32366) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1307) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5401) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28482) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26555) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7253) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20954) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9831) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26349) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12114) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4739) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29467) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9678) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26508) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11064) * $signed(input_fmap_33[7:0]) +
	( 11'sd 737) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_35[7:0]) +
	( 8'sd 114) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23938) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14763) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20941) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7501) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9171) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23617) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26594) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30950) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26051) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13682) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3440) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26865) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30553) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1667) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10224) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4978) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22886) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30595) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31965) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23149) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4972) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6024) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14430) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15587) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28251) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2226) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20508) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_87[7:0]) +
	( 11'sd 884) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3473) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32637) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4382) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28145) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28029) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13895) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29068) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8587) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8473) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2952) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9970) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14553) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4613) * $signed(input_fmap_109[7:0]) +
	( 10'sd 472) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14603) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26035) * $signed(input_fmap_112[7:0]) +
	( 10'sd 376) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7914) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8457) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10314) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29310) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20516) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14501) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 16'sd 24191) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21612) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32548) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26951) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27631) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8517) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13464) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13911) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4696) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5902) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2542) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17057) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11793) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2508) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28457) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5891) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1259) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2207) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_27[7:0]) +
	( 10'sd 354) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22229) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32086) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15098) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21329) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17366) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5405) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21947) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26790) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4344) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3518) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24700) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10421) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21878) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15256) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22718) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9977) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_54[7:0]) +
	( 10'sd 306) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23726) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6480) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24301) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2171) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28589) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6910) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16397) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9829) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26133) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13925) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17312) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31522) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23497) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18042) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24844) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23914) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20051) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11415) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7287) * $signed(input_fmap_90[7:0]) +
	( 10'sd 273) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28207) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31173) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11206) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29620) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22379) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12172) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6796) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23678) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15597) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2986) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24337) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8941) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7239) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23582) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12775) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7815) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27249) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22362) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18935) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 16'sd 22963) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19023) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9612) * $signed(input_fmap_2[7:0]) +
	( 11'sd 594) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26011) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11576) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25279) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11735) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23918) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9042) * $signed(input_fmap_10[7:0]) +
	( 14'sd 8163) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29847) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23294) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5152) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9625) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17700) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4328) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18669) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17683) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30838) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15146) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8890) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5265) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15605) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25737) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8707) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32410) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10522) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9261) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21969) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9199) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13325) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11510) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22803) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8625) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3561) * $signed(input_fmap_55[7:0]) +
	( 7'sd 56) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8608) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8390) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20107) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23441) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7606) * $signed(input_fmap_64[7:0]) +
	( 9'sd 207) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11440) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32014) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19947) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25944) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18250) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10675) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3742) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15724) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5895) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31420) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24612) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10528) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7801) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18765) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12257) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29888) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6701) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2692) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17178) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1638) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_102[7:0]) +
	( 7'sd 33) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6319) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26929) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18847) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31673) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4945) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9672) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21986) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1152) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3827) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16584) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16864) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_118[7:0]) +
	( 10'sd 333) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25847) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28049) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17916) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1664) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29863) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9296) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 14'sd 5472) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31959) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32060) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26867) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20670) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31146) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18693) * $signed(input_fmap_10[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9539) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24842) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25948) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4603) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8854) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14164) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27732) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20348) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3646) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6714) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13514) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24913) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31179) * $signed(input_fmap_27[7:0]) +
	( 11'sd 756) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3968) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11395) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2580) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16474) * $signed(input_fmap_37[7:0]) +
	( 8'sd 106) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4392) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17154) * $signed(input_fmap_40[7:0]) +
	( 10'sd 372) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6270) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25181) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28628) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3314) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16455) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22118) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27217) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14024) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19264) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16698) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1039) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32550) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11595) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19659) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13393) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6346) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9256) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16792) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14176) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6237) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29374) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25308) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_74[7:0]) +
	( 13'sd 4063) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10063) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4134) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13357) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6132) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10802) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10559) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13910) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6678) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22043) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29552) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26071) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26047) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31173) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21606) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16681) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17899) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9318) * $signed(input_fmap_100[7:0]) +
	( 11'sd 533) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14857) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7091) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28311) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29110) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19471) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1731) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26257) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29477) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30939) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26318) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28756) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1353) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15470) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21861) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1560) * $signed(input_fmap_124[7:0]) +
	( 11'sd 514) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8260) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 6'sd 27) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27264) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25474) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8917) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13617) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19511) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30746) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24220) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3573) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15037) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23502) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16466) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11404) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24435) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23535) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12779) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22987) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6123) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13630) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22326) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10925) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8901) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22774) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25174) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18879) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28324) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17764) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12028) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6536) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31508) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16408) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28817) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22649) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12654) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14252) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12349) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28755) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10488) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20549) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2249) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21181) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29332) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17663) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27213) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24046) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23736) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4683) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13152) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12446) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14847) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9105) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12658) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24269) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3220) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18363) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29198) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32613) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17698) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4666) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2290) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20509) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24570) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20742) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26550) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27260) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16879) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7088) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3043) * $signed(input_fmap_103[7:0]) +
	( 10'sd 266) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23083) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8438) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6243) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31366) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12683) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9926) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16761) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19203) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28537) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24999) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26000) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23529) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31061) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 16'sd 32288) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17589) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_2[7:0]) +
	( 10'sd 497) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17441) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10244) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24827) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23129) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24037) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25630) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18641) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16839) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16241) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17361) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27723) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24903) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27213) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4887) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31626) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8705) * $signed(input_fmap_26[7:0]) +
	( 10'sd 439) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20541) * $signed(input_fmap_28[7:0]) +
	( 11'sd 863) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28342) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26712) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17446) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26637) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4626) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2081) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31892) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32019) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11028) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26307) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32449) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8462) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16134) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1517) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29497) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2900) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14119) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8830) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13604) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28933) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4723) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6069) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_63[7:0]) +
	( 11'sd 519) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17691) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17595) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9167) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23123) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30844) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24742) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32180) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30203) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31569) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18643) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5674) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10669) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15614) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10244) * $signed(input_fmap_83[7:0]) +
	( 10'sd 454) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9635) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15208) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29317) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24939) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16927) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12519) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13888) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25061) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24495) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15279) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14575) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24289) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25466) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4221) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23963) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26147) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3761) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9258) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22957) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31926) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1768) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20243) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2764) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27836) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6965) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5103) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24842) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13740) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23967) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 16'sd 29276) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30552) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24879) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18334) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28125) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8172) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15054) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1278) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5231) * $signed(input_fmap_11[7:0]) +
	( 13'sd 4058) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22906) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26729) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4369) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20721) * $signed(input_fmap_19[7:0]) +
	( 7'sd 45) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15165) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5767) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24037) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16170) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3021) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4457) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16558) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3050) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22154) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20765) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25023) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10038) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17112) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27797) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7152) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10263) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16257) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27463) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8208) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7324) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5832) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23283) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6168) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1045) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28128) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3014) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18216) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3844) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5808) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2702) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9485) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21765) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27399) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10651) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30954) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23284) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23572) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7132) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14477) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1872) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29773) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28507) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_83[7:0]) +
	( 10'sd 284) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16354) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20722) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23045) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11173) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15047) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32441) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18139) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6575) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_95[7:0]) +
	( 11'sd 793) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9462) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24578) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2892) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18901) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19981) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32524) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11553) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1486) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21928) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28696) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23090) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23824) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24670) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13187) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 12'sd 1823) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17868) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23060) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1249) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4375) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18057) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24788) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22666) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21055) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8582) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1490) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24800) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28671) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13408) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28844) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15224) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28365) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10447) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26412) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5439) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14736) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24557) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12370) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25938) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18530) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30958) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26469) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25327) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12456) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23712) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21557) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6223) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5726) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3602) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32491) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19100) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30396) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6993) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10135) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1392) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6624) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24505) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19539) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22043) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11428) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10884) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13803) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14676) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10770) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30540) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10890) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17989) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4168) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7405) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22426) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1503) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31917) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18886) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31394) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6458) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6315) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24996) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10086) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27108) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9685) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17535) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25563) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1359) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19423) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29985) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3001) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20509) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1160) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18302) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18945) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29462) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18211) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24947) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27028) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 16'sd 22840) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23869) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5581) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7700) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18952) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30091) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28944) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7537) * $signed(input_fmap_12[7:0]) +
	( 11'sd 876) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10712) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17604) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29502) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28207) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20157) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30371) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19810) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_24[7:0]) +
	( 9'sd 158) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11927) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31512) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12761) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5567) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7210) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24365) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27730) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_34[7:0]) +
	( 12'sd 2007) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15657) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12200) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19409) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20256) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8356) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28452) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23195) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18954) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16074) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1737) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7815) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10401) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15643) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27560) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12745) * $signed(input_fmap_57[7:0]) +
	( 10'sd 395) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6154) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18766) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2292) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4510) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26901) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18115) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24207) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14863) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6237) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24847) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24940) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21220) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11300) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26355) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19705) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25409) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16588) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7035) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20570) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25336) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24817) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12192) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29569) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26350) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10948) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4822) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4742) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6191) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30978) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25323) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11903) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31101) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19472) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12975) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14925) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20857) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10360) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11066) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5411) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7145) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29536) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10491) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9786) * $signed(input_fmap_126[7:0]) +
	( 11'sd 793) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 15'sd 11229) * $signed(input_fmap_0[7:0]) +
	( 11'sd 974) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30737) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20828) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20149) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27970) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30175) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16201) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32750) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23486) * $signed(input_fmap_18[7:0]) +
	( 10'sd 350) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29581) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19721) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27066) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23340) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18849) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24971) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15578) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31507) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32476) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4476) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29713) * $signed(input_fmap_33[7:0]) +
	( 10'sd 498) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22069) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31503) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11527) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11174) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3613) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29054) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15204) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4725) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27791) * $signed(input_fmap_43[7:0]) +
	( 10'sd 435) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24226) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32738) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22583) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22153) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31764) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23214) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8218) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6277) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30272) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1920) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14195) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5589) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27614) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10508) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15773) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14376) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31123) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8045) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5131) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24649) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22784) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31779) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_78[7:0]) +
	( 9'sd 199) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20239) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20998) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15691) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21323) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11309) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32453) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20805) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6572) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1901) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2910) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26797) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5756) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30138) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_103[7:0]) +
	( 11'sd 997) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26179) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31068) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25104) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26341) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19219) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5551) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2152) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1774) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22367) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_118[7:0]) +
	( 11'sd 889) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8775) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23756) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2684) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1867) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6937) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 28810) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26031) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27262) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7265) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29080) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19164) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14363) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8517) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19940) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32535) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27916) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13538) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4968) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4871) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4702) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9624) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13905) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4890) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2093) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17781) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22628) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26303) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27293) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22614) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7294) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25119) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10985) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19407) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9515) * $signed(input_fmap_52[7:0]) +
	( 11'sd 1016) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22035) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8516) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13228) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16111) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9227) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27119) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18316) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11587) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21126) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7563) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13098) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22994) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24428) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3476) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6600) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8391) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6843) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8275) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18884) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15472) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28668) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26281) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25955) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18238) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3370) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12357) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9666) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12018) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22313) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3592) * $signed(input_fmap_93[7:0]) +
	( 11'sd 994) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12370) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22779) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29650) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18298) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23914) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20334) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5588) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8296) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1841) * $signed(input_fmap_107[7:0]) +
	( 11'sd 697) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23957) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6578) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20921) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13472) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21309) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2188) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31626) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15027) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10234) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 15'sd 10515) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7563) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18288) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19476) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12325) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11260) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13926) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21541) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6509) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3592) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32178) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3715) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21312) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13080) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29919) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26932) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21575) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6045) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17027) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20218) * $signed(input_fmap_29[7:0]) +
	( 4'sd 5) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13029) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24636) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18600) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28439) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18327) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15730) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19002) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25666) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26155) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18527) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26572) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_48[7:0]) +
	( 10'sd 508) * $signed(input_fmap_49[7:0]) +
	( 11'sd 795) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26941) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32532) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25122) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17061) * $signed(input_fmap_55[7:0]) +
	( 8'sd 113) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25416) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12964) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10306) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2744) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31796) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19627) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6283) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22800) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7560) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14619) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25372) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31976) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1030) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7963) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12744) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18080) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29020) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7840) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24932) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28333) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10457) * $signed(input_fmap_84[7:0]) +
	( 11'sd 987) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19095) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15311) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18760) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29023) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12518) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14084) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20779) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21373) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6285) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9436) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5375) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6324) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6250) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18250) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28681) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3254) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20432) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27241) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19140) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9226) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13324) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23084) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17735) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3799) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 15'sd 14343) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29800) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8540) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21022) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_4[7:0]) +
	( 11'sd 582) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1668) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_7[7:0]) +
	( 11'sd 1021) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12724) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29198) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2831) * $signed(input_fmap_11[7:0]) +
	( 10'sd 383) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15476) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23175) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26524) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18348) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4555) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11361) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28483) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14182) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16827) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13503) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19797) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_27[7:0]) +
	( 9'sd 250) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12248) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5588) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5475) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18769) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31663) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4526) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_40[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_41[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31500) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17015) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4383) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6892) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32498) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17955) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26526) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26050) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32697) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3484) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3337) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12729) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22511) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23628) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28382) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12810) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26271) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32537) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4617) * $signed(input_fmap_75[7:0]) +
	( 11'sd 989) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26844) * $signed(input_fmap_77[7:0]) +
	( 7'sd 53) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7523) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28668) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8529) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5138) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25890) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20450) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20434) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17114) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29880) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20396) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18330) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4627) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12014) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5105) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1815) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17563) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5767) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13800) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14689) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31963) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31718) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7905) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28924) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19966) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28976) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10860) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9837) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29943) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31330) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11759) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16478) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11538) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20636) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20842) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4900) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26860) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11968) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 16'sd 16714) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6570) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7744) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2489) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4418) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21703) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6000) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6100) * $signed(input_fmap_9[7:0]) +
	( 11'sd 664) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30686) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26120) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17160) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25809) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18898) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22101) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30351) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19615) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29199) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14347) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4450) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22294) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24282) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25491) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15111) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1154) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3968) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5410) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16149) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8883) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32390) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13704) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18688) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21784) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19783) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25537) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15376) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14985) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12654) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13537) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11363) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26183) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15731) * $signed(input_fmap_66[7:0]) +
	( 11'sd 896) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19478) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3780) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8112) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19044) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28758) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27726) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20387) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4100) * $signed(input_fmap_78[7:0]) +
	( 11'sd 962) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4404) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30905) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31569) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8220) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15499) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31539) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3234) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23510) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8918) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20192) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14283) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23912) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17910) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32716) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20493) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7050) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8820) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31779) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11222) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10622) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14246) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19327) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14636) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24622) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17527) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6504) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15310) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4167) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17192) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2810) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 16'sd 24076) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27801) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_2[7:0]) +
	( 8'sd 119) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10693) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11421) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16525) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31083) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22353) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15905) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14658) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6493) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15183) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6972) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32097) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30311) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5793) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30422) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25355) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6665) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21133) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_30[7:0]) +
	( 9'sd 177) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_32[7:0]) +
	( 10'sd 353) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32147) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22926) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6803) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5807) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18828) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27941) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4430) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19615) * $signed(input_fmap_46[7:0]) +
	( 10'sd 482) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8974) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29148) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11330) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13308) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16622) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21093) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29759) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14147) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23501) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25906) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8846) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17245) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20047) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30897) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28442) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1463) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21767) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20471) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18030) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3918) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8780) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9661) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16845) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16573) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8741) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27563) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7732) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31480) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28164) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21461) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12972) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31173) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22636) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1680) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30127) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_97[7:0]) +
	( 4'sd 4) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16946) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1390) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30567) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3713) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7943) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21480) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31340) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7749) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28367) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1991) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14473) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24713) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16489) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4270) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 16'sd 20216) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7747) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11855) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31304) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32116) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17670) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9691) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_10[7:0]) +
	( 11'sd 858) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6980) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11036) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29776) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28819) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3875) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16627) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22617) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32167) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26933) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1418) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13686) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2243) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22263) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2749) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6905) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32681) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8730) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8783) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11173) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7578) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14776) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12966) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7433) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3068) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13164) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3870) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14885) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4715) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26016) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5359) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7777) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22238) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20783) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22914) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21685) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4271) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19001) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31724) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4818) * $signed(input_fmap_81[7:0]) +
	( 8'sd 65) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1866) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28797) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21312) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4375) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14019) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13547) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12268) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31687) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13878) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31806) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20153) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16483) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13977) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22239) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10147) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29065) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12504) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24865) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30780) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16497) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16896) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4867) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1870) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28141) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5927) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2305) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8828) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30278) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30309) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 14'sd 6971) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28873) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30969) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15912) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5041) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1900) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12104) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23326) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31298) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32761) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9594) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14361) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13242) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18917) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4328) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6854) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11449) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23100) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25651) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10365) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2353) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24243) * $signed(input_fmap_37[7:0]) +
	( 11'sd 938) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21512) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16182) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29503) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23072) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2644) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25415) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11820) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11699) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17880) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6896) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24903) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13931) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14444) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8156) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16388) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30054) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13788) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16262) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_64[7:0]) +
	( 11'sd 813) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5495) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27338) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32360) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12831) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22303) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21395) * $signed(input_fmap_77[7:0]) +
	( 11'sd 553) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_81[7:0]) +
	( 9'sd 175) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14792) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15592) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7343) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3492) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25563) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27177) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7470) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15851) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26944) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5020) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25254) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27315) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4642) * $signed(input_fmap_102[7:0]) +
	( 10'sd 495) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13679) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2318) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4755) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12925) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5804) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_111[7:0]) +
	( 11'sd 665) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11359) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32242) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9827) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5027) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22676) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8279) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8370) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9998) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10294) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25315) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10953) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24277) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 16'sd 22831) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24177) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3626) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20532) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9191) * $signed(input_fmap_4[7:0]) +
	( 10'sd 477) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19370) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28696) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23584) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11640) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19265) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6538) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28311) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28265) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3206) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30281) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23463) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18496) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29898) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6247) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11327) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31986) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29923) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24776) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29829) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20595) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5815) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7741) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14617) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8337) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23996) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10334) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7704) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9569) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18125) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1347) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19612) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23576) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1640) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32574) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31905) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28032) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1797) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28115) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4129) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22374) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9105) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2239) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29289) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13292) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12416) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7795) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18420) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3689) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13271) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22404) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28511) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19251) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7986) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21644) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10003) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16301) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30448) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16008) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12410) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27891) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19253) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22347) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19616) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19618) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4498) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29980) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31180) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2990) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2744) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27517) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27119) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13056) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26622) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26678) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11797) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6556) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24935) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 15'sd 11793) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11795) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9610) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28929) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11531) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1877) * $signed(input_fmap_6[7:0]) +
	( 11'sd 689) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17250) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14873) * $signed(input_fmap_9[7:0]) +
	( 10'sd 348) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31233) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20081) * $signed(input_fmap_14[7:0]) +
	( 10'sd 426) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13537) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27216) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4302) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29465) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12324) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27022) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5703) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2155) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4991) * $signed(input_fmap_29[7:0]) +
	( 12'sd 2010) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28558) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30969) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26752) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23054) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2268) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_41[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14275) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4259) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26470) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31427) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_49[7:0]) +
	( 9'sd 132) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19160) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22076) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24354) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6042) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19260) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23395) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28476) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26955) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27072) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26791) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12960) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6998) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23923) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_69[7:0]) +
	( 11'sd 597) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29195) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30863) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16350) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25605) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13608) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13279) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30127) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6716) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27938) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11719) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25776) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2737) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27514) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32446) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11183) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10714) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31985) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9877) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22497) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28236) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4984) * $signed(input_fmap_108[7:0]) +
	( 10'sd 375) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17304) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13689) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11706) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28103) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32295) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5696) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24721) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17215) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 12'sd 1399) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2075) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31986) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15781) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21681) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28177) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15009) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5999) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30085) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9017) * $signed(input_fmap_14[7:0]) +
	( 9'sd 192) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11152) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5248) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2153) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15692) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10978) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4514) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27784) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28267) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6905) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22467) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7241) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30111) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16974) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3928) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22300) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10401) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14919) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1095) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6325) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1664) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15622) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18819) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13777) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31843) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8692) * $signed(input_fmap_58[7:0]) +
	( 8'sd 74) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5709) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29675) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7421) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25296) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29397) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23350) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12643) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7869) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_73[7:0]) +
	( 10'sd 350) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20350) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31582) * $signed(input_fmap_76[7:0]) +
	( 10'sd 300) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30264) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29794) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6532) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10685) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1501) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14402) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24606) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10338) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32052) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27304) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21744) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9206) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8609) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8200) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30521) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13248) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27916) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19986) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_104[7:0]) +
	( 11'sd 662) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30045) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7561) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18400) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14283) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_113[7:0]) +
	( 11'sd 700) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10870) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1353) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11775) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16887) * $signed(input_fmap_120[7:0]) +
	( 11'sd 641) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10793) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23182) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11355) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18218) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32199) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 14'sd 6599) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7337) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2710) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8248) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6818) * $signed(input_fmap_4[7:0]) +
	( 10'sd 456) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3370) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23771) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4401) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22325) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19431) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15228) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15313) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26323) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28939) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6913) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4239) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24861) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6512) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30883) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32684) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24431) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26876) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8591) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27330) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2702) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15806) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28176) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20269) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_48[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6219) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5311) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11690) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31105) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28358) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10381) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30363) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5513) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20895) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3723) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18213) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13575) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17091) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3467) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16158) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25630) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_68[7:0]) +
	( 10'sd 510) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10437) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11738) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2357) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22025) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30242) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29896) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7319) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1725) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11004) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23496) * $signed(input_fmap_81[7:0]) +
	( 11'sd 785) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14682) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18487) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25292) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6470) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24035) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17837) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5490) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2326) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10189) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26725) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16913) * $signed(input_fmap_95[7:0]) +
	( 14'sd 8090) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28721) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22902) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5059) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5236) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21991) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4763) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31379) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11961) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9636) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29643) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1983) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27184) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16590) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14606) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6848) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20704) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29993) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10116) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25544) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23058) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 15'sd 11616) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1907) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10705) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14730) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20881) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10348) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8616) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29305) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10556) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30463) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28922) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4426) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9893) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13768) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29436) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19163) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20013) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8052) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3331) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6879) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21860) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8234) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27091) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30321) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9017) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5464) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10222) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32421) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1422) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29663) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8310) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18602) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22802) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12360) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1160) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6107) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22373) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30899) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22995) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12468) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6606) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18703) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28033) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9761) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11573) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10931) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21909) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23409) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_77[7:0]) +
	( 9'sd 226) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29169) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2094) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_82[7:0]) +
	( 13'sd 4027) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31625) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30426) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12739) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11671) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_92[7:0]) +
	( 11'sd 704) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22303) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2980) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6230) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20434) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13907) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31105) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13610) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20609) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23558) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5011) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6156) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27072) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12503) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31130) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1552) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11445) * $signed(input_fmap_116[7:0]) +
	( 9'sd 231) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4190) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16822) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23684) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15430) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5868) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20608) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 15'sd 16147) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16606) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9316) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1228) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29653) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29955) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28833) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31815) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25857) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22599) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4941) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22445) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28885) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23668) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1618) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21244) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15761) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15218) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4554) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4212) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7424) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32735) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15702) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15474) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16194) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_33[7:0]) +
	( 10'sd 468) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5252) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3603) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25404) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18155) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21803) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24597) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19869) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18256) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22118) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23047) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20194) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29116) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22930) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26837) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31382) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18955) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8876) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12154) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31575) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15753) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30046) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4721) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20274) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23728) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7518) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26021) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12745) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24020) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5550) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23169) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22024) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30856) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5854) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19938) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21588) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7422) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23999) * $signed(input_fmap_96[7:0]) +
	( 11'sd 554) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18382) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14459) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22259) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16871) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20768) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28270) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25150) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5970) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3658) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31584) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20818) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20717) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11420) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23434) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14891) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14419) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4170) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11503) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6084) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25431) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20129) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4657) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24184) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 16'sd 30746) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12985) * $signed(input_fmap_1[7:0]) +
	( 10'sd 434) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28524) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8088) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17998) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28079) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7403) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24061) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14393) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3449) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2555) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4621) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9212) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3895) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3175) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9568) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28471) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18363) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27105) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31305) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18274) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21318) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7729) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4021) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20802) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29260) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14263) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_38[7:0]) +
	( 10'sd 477) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24132) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14652) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7484) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6315) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10567) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12799) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19294) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17430) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19368) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26384) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16122) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12507) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24406) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29976) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18081) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15429) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30739) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26964) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27658) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26730) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26530) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19728) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31682) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16230) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21006) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12751) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26331) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5155) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16854) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28913) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5207) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13093) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13095) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31975) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11973) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30777) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26193) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20977) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28666) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16422) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1604) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9644) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5627) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1034) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12177) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5659) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16682) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26192) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18894) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28828) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8173) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1216) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6512) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21783) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29669) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5383) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30135) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_125[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27947) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 14'sd 4898) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17209) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32506) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16330) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15163) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18959) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23250) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25894) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14473) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31944) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5316) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5555) * $signed(input_fmap_15[7:0]) +
	( 10'sd 389) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15318) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16691) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7530) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25513) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26136) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1699) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14804) * $signed(input_fmap_24[7:0]) +
	( 10'sd 305) * $signed(input_fmap_25[7:0]) +
	( 9'sd 212) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28536) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7014) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28537) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6364) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26211) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21485) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4044) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28082) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17230) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22040) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26348) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26036) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29234) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7644) * $signed(input_fmap_46[7:0]) +
	( 11'sd 773) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10850) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14286) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2361) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1823) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14311) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25591) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25732) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10270) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5452) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23039) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25651) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_68[7:0]) +
	( 9'sd 250) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11769) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25239) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12510) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22332) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13782) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8510) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30682) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30631) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13112) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16299) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10814) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26016) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14508) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13325) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24957) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12142) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15679) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3977) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31460) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7989) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7666) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27569) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6917) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29713) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4829) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3967) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3799) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21334) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17550) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27826) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29350) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23730) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2511) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31754) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32535) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 16'sd 25185) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21919) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30967) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31897) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5021) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23093) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4946) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24856) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2528) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21175) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8573) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1934) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_20[7:0]) +
	( 13'sd 4076) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15285) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5796) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30001) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27034) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23751) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26779) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32048) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1832) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11633) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24020) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27983) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18247) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21772) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18867) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3227) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27568) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1349) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2183) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29756) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22864) * $signed(input_fmap_50[7:0]) +
	( 10'sd 431) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18752) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25491) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25882) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17096) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13598) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17970) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21936) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15210) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16843) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22217) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6887) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4397) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12920) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_75[7:0]) +
	( 10'sd 319) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31039) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23063) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14948) * $signed(input_fmap_84[7:0]) +
	( 13'sd 4007) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31578) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28174) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18556) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12346) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32692) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4734) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_97[7:0]) +
	( 14'sd 8127) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14125) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13380) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15733) * $signed(input_fmap_103[7:0]) +
	( 6'sd 27) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8402) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6457) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23288) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24218) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19774) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28476) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24558) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8521) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5739) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26736) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14402) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28730) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24509) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11951) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12007) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2578) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28645) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 16'sd 30144) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8621) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3253) * $signed(input_fmap_3[7:0]) +
	( 11'sd 919) * $signed(input_fmap_4[7:0]) +
	( 11'sd 902) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28489) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18228) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21337) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2264) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28272) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7948) * $signed(input_fmap_14[7:0]) +
	( 10'sd 400) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12150) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10191) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28019) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30323) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27408) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8582) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19692) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21774) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26791) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7739) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4337) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10760) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31981) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3484) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1858) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10055) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6202) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9913) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3708) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2685) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6129) * $signed(input_fmap_47[7:0]) +
	( 11'sd 841) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15451) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24861) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28984) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16556) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5111) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1902) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32450) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14976) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23953) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17427) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30661) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11598) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28151) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26473) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27924) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27269) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20879) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22480) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26363) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9037) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32118) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19127) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19794) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20822) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25248) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24460) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14703) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21319) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30495) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6201) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14795) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22095) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31412) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5177) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13913) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19632) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6723) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9220) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9183) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5218) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15413) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 16'sd 21600) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4898) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7330) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29464) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_6[7:0]) +
	( 11'sd 917) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26537) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32581) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4500) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10864) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13689) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16072) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4484) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_19[7:0]) +
	( 11'sd 933) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32492) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_25[7:0]) +
	( 9'sd 188) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20683) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12924) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11234) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9830) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31281) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3206) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31539) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11166) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32328) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31499) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19768) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7466) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11892) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3280) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24693) * $signed(input_fmap_49[7:0]) +
	( 9'sd 170) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8429) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8840) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2681) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9031) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20843) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14509) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9019) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14784) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_66[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_71[7:0]) +
	( 10'sd 338) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28793) * $signed(input_fmap_73[7:0]) +
	( 11'sd 724) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27770) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17044) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26059) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8294) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13099) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3115) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31567) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6044) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6611) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29304) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30127) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24892) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14220) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19879) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14026) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10759) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21765) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18738) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8698) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18795) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5368) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29664) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13158) * $signed(input_fmap_110[7:0]) +
	( 10'sd 450) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12796) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18290) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9096) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18678) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11368) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1492) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17647) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6605) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4459) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21489) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9549) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22952) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 16'sd 30070) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16283) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16064) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27887) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27992) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31944) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13833) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19012) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11666) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15687) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31837) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9651) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19420) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17142) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19508) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4565) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10050) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30076) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14224) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8640) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17331) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15208) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19054) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30542) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20774) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28910) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20764) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11018) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2652) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12167) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28604) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7766) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31912) * $signed(input_fmap_53[7:0]) +
	( 6'sd 18) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15870) * $signed(input_fmap_55[7:0]) +
	( 9'sd 135) * $signed(input_fmap_56[7:0]) +
	( 11'sd 554) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13094) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13020) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30004) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10402) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8376) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19773) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25982) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14632) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7876) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11765) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15941) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26640) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21701) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16498) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24113) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18006) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8470) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2798) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11537) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31218) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15068) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18530) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29779) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7640) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13311) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4718) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19509) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26977) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2692) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9350) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24728) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1223) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15410) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24242) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23550) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6874) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6540) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25084) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6357) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28309) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22572) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1130) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11025) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17989) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17165) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 15'sd 15178) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13265) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8209) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23741) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1900) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_5[7:0]) +
	( 10'sd 396) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21146) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13519) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28089) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4305) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3218) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15634) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1476) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15553) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30048) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19650) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24570) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4347) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22266) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13888) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19056) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22669) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11505) * $signed(input_fmap_31[7:0]) +
	( 11'sd 897) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5465) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17867) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30255) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26279) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29728) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7023) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17979) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30600) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18013) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14877) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13177) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18988) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20981) * $signed(input_fmap_45[7:0]) +
	( 11'sd 753) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8111) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14360) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27013) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24151) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_52[7:0]) +
	( 11'sd 617) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1526) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30052) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5959) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12686) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26549) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28150) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27222) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25225) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23134) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23315) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5903) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22616) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13007) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31815) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25508) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2878) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13013) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25038) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29065) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10713) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17649) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11974) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11697) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9708) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8535) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5610) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10927) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22803) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5597) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1392) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8205) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20012) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24124) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2669) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15181) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15632) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16569) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31787) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15761) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25368) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6806) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13009) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3474) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24130) * $signed(input_fmap_115[7:0]) +
	( 10'sd 388) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29087) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10414) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6937) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26599) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_122[7:0]) +
	( 11'sd 853) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 14'sd 6509) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15938) * $signed(input_fmap_1[7:0]) +
	( 11'sd 905) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14718) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14678) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30253) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27341) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8348) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31832) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26752) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11480) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12014) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1516) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28983) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12418) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18611) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17851) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12795) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17062) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22317) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19215) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6932) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25242) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31320) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8492) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4215) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14115) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3897) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7718) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29291) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22009) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31345) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6180) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31804) * $signed(input_fmap_46[7:0]) +
	( 10'sd 468) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4797) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26749) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19452) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15650) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3180) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15010) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28333) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20588) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1782) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24850) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4191) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24165) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18552) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5904) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3177) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2635) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3459) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15087) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17058) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17098) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15652) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30238) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13090) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2117) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7328) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_87[7:0]) +
	( 11'sd 1022) * $signed(input_fmap_88[7:0]) +
	( 10'sd 387) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8642) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18686) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26448) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6026) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13886) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20678) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11912) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9451) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27692) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16617) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6727) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14223) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18323) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20192) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31132) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18690) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16643) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_117[7:0]) +
	( 10'sd 448) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9209) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20339) * $signed(input_fmap_122[7:0]) +
	( 11'sd 749) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3135) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25620) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 13'sd 2640) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2191) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28488) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19762) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11492) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20750) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5959) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32004) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32699) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19795) * $signed(input_fmap_14[7:0]) +
	( 10'sd 464) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22687) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24039) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29065) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30948) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26464) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5123) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13280) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21879) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13447) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10385) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25057) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12064) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11678) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31396) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26570) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25815) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16401) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30450) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6616) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17129) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12378) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22087) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23143) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19827) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23382) * $signed(input_fmap_51[7:0]) +
	( 10'sd 483) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14724) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16482) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28983) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4239) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7049) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4120) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25649) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24106) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_64[7:0]) +
	( 11'sd 586) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14428) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2296) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10865) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28111) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24713) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1585) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9349) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6951) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19994) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9173) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10499) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30615) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16623) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26190) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13102) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9865) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23558) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13694) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14578) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27654) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29304) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7080) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29214) * $signed(input_fmap_101[7:0]) +
	( 8'sd 67) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4471) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30493) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24194) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7213) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25598) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6172) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6849) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25645) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2764) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23537) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17356) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24512) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 16'sd 22624) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21114) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3081) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24696) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30476) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30406) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18618) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20791) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7661) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29334) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17201) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21412) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_20[7:0]) +
	( 8'sd 127) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26766) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18243) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24349) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12849) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2965) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9524) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23867) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15465) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20966) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19560) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31600) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4726) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22215) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32119) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31961) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27376) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12333) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17347) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5822) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24736) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9352) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10449) * $signed(input_fmap_58[7:0]) +
	( 10'sd 307) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20282) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28123) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25098) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3478) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11081) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17678) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22302) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31956) * $signed(input_fmap_71[7:0]) +
	( 13'sd 4009) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17044) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5056) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19655) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27958) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29110) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32081) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19483) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27624) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29860) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1538) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10412) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18146) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28118) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21417) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24599) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26912) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26002) * $signed(input_fmap_103[7:0]) +
	( 12'sd 2039) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8528) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7025) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31211) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15877) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21099) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4571) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13105) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25995) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20137) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1991) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25202) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15379) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32204) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25050) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17366) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 16'sd 30880) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5907) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1093) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22804) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21763) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1503) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11069) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1926) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9387) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29270) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20492) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23023) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26921) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17618) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29441) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24479) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23847) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20754) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25829) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21926) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8507) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1488) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30833) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_37[7:0]) +
	( 11'sd 619) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1892) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19814) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29222) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23639) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25258) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5458) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29943) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8201) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21362) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32401) * $signed(input_fmap_65[7:0]) +
	( 9'sd 214) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14737) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16445) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14119) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21750) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18782) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6409) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_78[7:0]) +
	( 10'sd 389) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24216) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30489) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31450) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6113) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18858) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21059) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32542) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16554) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29533) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13002) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29752) * $signed(input_fmap_97[7:0]) +
	( 11'sd 656) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26709) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6408) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18795) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21237) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31801) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16181) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8176) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12449) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26873) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25177) * $signed(input_fmap_114[7:0]) +
	( 11'sd 785) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13905) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_117[7:0]) +
	( 9'sd 132) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22778) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14453) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1691) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 14'sd 7603) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30948) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22174) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13610) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10689) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1714) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19569) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12181) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1966) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4514) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6634) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10712) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_16[7:0]) +
	( 13'sd 4067) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10876) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18490) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23617) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15888) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23301) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8328) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5513) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5483) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22140) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6524) * $signed(input_fmap_34[7:0]) +
	( 11'sd 735) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5322) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1772) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21017) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27510) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27080) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20498) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23736) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21839) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10840) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26776) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5905) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15062) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11207) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17590) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17566) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20178) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23902) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21687) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19867) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14031) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14194) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9496) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_71[7:0]) +
	( 7'sd 53) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15363) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21841) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14493) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28907) * $signed(input_fmap_78[7:0]) +
	( 9'sd 154) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9681) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11215) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27640) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29439) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15915) * $signed(input_fmap_89[7:0]) +
	( 11'sd 950) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15706) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12090) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26810) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21517) * $signed(input_fmap_97[7:0]) +
	( 14'sd 8073) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10076) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23964) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32720) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25465) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6963) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16442) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19855) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2638) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24989) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10416) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24468) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_120[7:0]) +
	( 9'sd 244) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28961) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4902) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12950) * $signed(input_fmap_126[7:0]) +
	( 11'sd 955) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 15'sd 14205) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29866) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1437) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_4[7:0]) +
	( 7'sd 48) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15380) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23921) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16525) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28791) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30153) * $signed(input_fmap_13[7:0]) +
	( 9'sd 186) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17902) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28183) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31222) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11959) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4144) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12892) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16920) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28793) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19589) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14337) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9116) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12299) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21397) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16344) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1556) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22931) * $signed(input_fmap_39[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19802) * $signed(input_fmap_41[7:0]) +
	( 12'sd 2031) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3571) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31708) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12942) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3628) * $signed(input_fmap_49[7:0]) +
	( 10'sd 352) * $signed(input_fmap_50[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8130) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7152) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29524) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15954) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26090) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4565) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15055) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5422) * $signed(input_fmap_68[7:0]) +
	( 10'sd 340) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13081) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24771) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28371) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3134) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12990) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32756) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22930) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6243) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29993) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22269) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32649) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3361) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29493) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21088) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17409) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9108) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30052) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13067) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2643) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29158) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29351) * $signed(input_fmap_103[7:0]) +
	( 11'sd 885) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7456) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24293) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15887) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9549) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4985) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21085) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4326) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1357) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28549) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26679) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5580) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16251) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22721) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7271) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22977) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 13'sd 3697) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32212) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20500) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12560) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11621) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5499) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6284) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29464) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17073) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32491) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22159) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19039) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13524) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9211) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32256) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26394) * $signed(input_fmap_17[7:0]) +
	( 13'sd 4048) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9672) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29642) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11001) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_22[7:0]) +
	( 13'sd 4009) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31372) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16986) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25351) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30640) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28835) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17433) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27329) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7203) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10437) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13855) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13762) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16175) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31662) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8651) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16020) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25525) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2285) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12797) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11800) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12995) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3637) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23167) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20532) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11094) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21650) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12073) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11126) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15953) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20000) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23910) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20089) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10093) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17612) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31604) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8566) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17775) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2562) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29965) * $signed(input_fmap_77[7:0]) +
	( 13'sd 4084) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10788) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10208) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12604) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31973) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11756) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30865) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13057) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15114) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25821) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30079) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21099) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3907) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21464) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9343) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2091) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24916) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29927) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18866) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9999) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14102) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31682) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13201) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15406) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_116[7:0]) +
	( 12'sd 2033) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_118[7:0]) +
	( 11'sd 561) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4785) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6846) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19282) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23885) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 14'sd 7526) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3915) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18846) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3737) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30126) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29682) * $signed(input_fmap_6[7:0]) +
	( 9'sd 142) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27260) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1037) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19723) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15761) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25883) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7704) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15408) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9999) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18951) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32675) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22004) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5318) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24934) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16081) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24116) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31359) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13205) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18869) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17412) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10773) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24976) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5999) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24138) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8669) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18163) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25105) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22512) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2637) * $signed(input_fmap_47[7:0]) +
	( 11'sd 512) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32453) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4906) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29956) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8223) * $signed(input_fmap_52[7:0]) +
	( 11'sd 553) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4589) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23698) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14290) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20509) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1130) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25820) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14918) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6061) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19065) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5418) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22727) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32085) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30641) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31102) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11365) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15600) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26280) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30723) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19407) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26433) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28462) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16215) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24180) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3490) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12666) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13039) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3416) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32374) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31452) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11425) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22606) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17801) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20961) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18506) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17772) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21004) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24721) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17517) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_111[7:0]) +
	( 10'sd 430) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15382) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18126) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29686) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22131) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1869) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1438) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19921) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9584) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 16'sd 16635) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3328) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25826) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5927) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32283) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8764) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10264) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19223) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16002) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13072) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12272) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5109) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17224) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16977) * $signed(input_fmap_23[7:0]) +
	( 11'sd 561) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4629) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4856) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26897) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8847) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1710) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31621) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25246) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29130) * $signed(input_fmap_38[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31435) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21204) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4731) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20397) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24770) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6262) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5559) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10283) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22238) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21802) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1039) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27423) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21807) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8588) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7289) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16756) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2539) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17156) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28277) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2715) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17333) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17695) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9688) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7849) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9660) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21838) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26874) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10161) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6727) * $signed(input_fmap_86[7:0]) +
	( 14'sd 8127) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8229) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23199) * $signed(input_fmap_90[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2937) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26367) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4329) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12485) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3970) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27850) * $signed(input_fmap_100[7:0]) +
	( 10'sd 406) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27517) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14366) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10612) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19792) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25636) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5976) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9661) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21590) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27497) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3072) * $signed(input_fmap_117[7:0]) +
	( 11'sd 1022) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8497) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18362) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18469) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4852) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16745) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14171) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 11'sd 955) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22610) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14658) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29868) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27605) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28539) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25531) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12296) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3645) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7061) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15505) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_15[7:0]) +
	( 11'sd 777) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30981) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12034) * $signed(input_fmap_18[7:0]) +
	( 10'sd 259) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24265) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23013) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9542) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27735) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5464) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4208) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9203) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12651) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14529) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18922) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18174) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2379) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19140) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17842) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4945) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14301) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12570) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13414) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29631) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32708) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5931) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6995) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30465) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7016) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17428) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14566) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32384) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27594) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8892) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10164) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8457) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18741) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28330) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7611) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14366) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28553) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_84[7:0]) +
	( 11'sd 870) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27070) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19462) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30251) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17122) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4479) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21994) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3557) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_100[7:0]) +
	( 14'sd 8059) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29212) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1279) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9501) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2810) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17133) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25781) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5331) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28993) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28973) * $signed(input_fmap_117[7:0]) +
	( 9'sd 226) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19152) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5557) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23160) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31683) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31047) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30334) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 15'sd 12800) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17612) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_4[7:0]) +
	( 10'sd 423) * $signed(input_fmap_5[7:0]) +
	( 9'sd 144) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1543) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22717) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3686) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4916) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17937) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25198) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1050) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29689) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31302) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3792) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6951) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15394) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31973) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11388) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2603) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2113) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3411) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28990) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1912) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12871) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_39[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21760) * $signed(input_fmap_45[7:0]) +
	( 14'sd 8055) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_47[7:0]) +
	( 14'sd 8001) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21924) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16478) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1238) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4611) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11172) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28084) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6019) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20995) * $signed(input_fmap_65[7:0]) +
	( 10'sd 331) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13688) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2602) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22724) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31910) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11140) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2325) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4543) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29317) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32453) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22609) * $signed(input_fmap_76[7:0]) +
	( 11'sd 584) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1370) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10075) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7439) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21624) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4699) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12846) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18648) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_91[7:0]) +
	( 5'sd 9) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_95[7:0]) +
	( 11'sd 863) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3732) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4358) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29222) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6222) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25628) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3301) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4984) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32001) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19289) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7926) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13935) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21379) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9006) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28760) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 16'sd 27195) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20317) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8224) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14864) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2133) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7238) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2304) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29061) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18006) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9139) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25269) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22316) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31365) * $signed(input_fmap_19[7:0]) +
	( 9'sd 252) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7530) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1602) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15092) * $signed(input_fmap_30[7:0]) +
	( 12'sd 2010) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5141) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2540) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14759) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13482) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21212) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26296) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32430) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3470) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23314) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15596) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9572) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16136) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2257) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10459) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19415) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17597) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8240) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26206) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15753) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21007) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16449) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5481) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2781) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25936) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11642) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8763) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4712) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29279) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15812) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25732) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18776) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26269) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22778) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6893) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10248) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10111) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9542) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7187) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4098) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29449) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26111) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30419) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1590) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26932) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27733) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19597) * $signed(input_fmap_104[7:0]) +
	( 9'sd 210) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26142) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16402) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3548) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14628) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13268) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27797) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9432) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13020) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21096) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12850) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5776) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 15'sd 9291) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24859) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7085) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7276) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7964) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1914) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25738) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9990) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27306) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9090) * $signed(input_fmap_13[7:0]) +
	( 10'sd 350) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8228) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_17[7:0]) +
	( 13'sd 4024) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31170) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20655) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20509) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9759) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9787) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24592) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17802) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4521) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16115) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11603) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_35[7:0]) +
	( 9'sd 231) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12460) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4946) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_42[7:0]) +
	( 10'sd 340) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24523) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5062) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13989) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11254) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4209) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9486) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28870) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9038) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28708) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5459) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28269) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10053) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13816) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16934) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31832) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3783) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27187) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15384) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12744) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5476) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23258) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8807) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21483) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25150) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8688) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23736) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16288) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8762) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23329) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_90[7:0]) +
	( 9'sd 130) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12948) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4301) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5054) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31522) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32705) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4169) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7215) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6887) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16418) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23342) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22593) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20600) * $signed(input_fmap_111[7:0]) +
	( 9'sd 164) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13398) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30068) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4878) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23935) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_120[7:0]) +
	( 10'sd 257) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17093) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17433) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21732) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31004) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 16'sd 22287) * $signed(input_fmap_0[7:0]) +
	( 8'sd 92) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19781) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22607) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5739) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7613) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29820) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27642) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30363) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20608) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23009) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18791) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25019) * $signed(input_fmap_18[7:0]) +
	( 11'sd 1010) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23794) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32069) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17314) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28049) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6788) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29033) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12969) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14166) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28924) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13022) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_33[7:0]) +
	( 8'sd 71) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15326) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31738) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19443) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4286) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18615) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4405) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8291) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22008) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20001) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12882) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23421) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_58[7:0]) +
	( 11'sd 534) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1452) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17477) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5441) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6225) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12615) * $signed(input_fmap_69[7:0]) +
	( 7'sd 56) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31010) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30511) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17770) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24159) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19090) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25213) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23115) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14293) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_84[7:0]) +
	( 10'sd 481) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20503) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20328) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31783) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21011) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10583) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16806) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21818) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2666) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1426) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7811) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4333) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16270) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21707) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7092) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7042) * $signed(input_fmap_106[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31881) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18518) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24027) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2171) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23694) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5996) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15975) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25920) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12377) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25050) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 16'sd 20535) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16135) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7067) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25770) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30917) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23518) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5299) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18894) * $signed(input_fmap_10[7:0]) +
	( 13'sd 4060) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9102) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11167) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13245) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15735) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29591) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5594) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25203) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9931) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17042) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_32[7:0]) +
	( 10'sd 338) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1908) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3101) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11843) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20765) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13653) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15772) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_46[7:0]) +
	( 10'sd 494) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28866) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14817) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4629) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15865) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28557) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23649) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31300) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27923) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22330) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15618) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12672) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12344) * $signed(input_fmap_66[7:0]) +
	( 9'sd 248) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31670) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3468) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21953) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27775) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29169) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10133) * $signed(input_fmap_76[7:0]) +
	( 11'sd 966) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3470) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25096) * $signed(input_fmap_79[7:0]) +
	( 11'sd 947) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32671) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22839) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29942) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2122) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27490) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18028) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25285) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30921) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23874) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3138) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23400) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6466) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11338) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19676) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4413) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31017) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23221) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_102[7:0]) +
	( 9'sd 223) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3010) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23403) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8857) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13206) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21699) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8498) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1467) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32096) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2757) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20070) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3932) * $signed(input_fmap_123[7:0]) +
	( 14'sd 8013) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10465) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6566) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 10'sd 296) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19853) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18128) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22850) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6302) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4636) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15127) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18775) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12729) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9405) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23366) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22249) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7697) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2149) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22102) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17354) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19873) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31140) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10319) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4111) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12200) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7382) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5430) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20962) * $signed(input_fmap_33[7:0]) +
	( 11'sd 790) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20136) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18458) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12274) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6148) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14270) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25266) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18999) * $signed(input_fmap_43[7:0]) +
	( 12'sd 2030) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24662) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3016) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26139) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7754) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31969) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11648) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7824) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5713) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_63[7:0]) +
	( 11'sd 847) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4937) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6983) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8352) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15445) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23596) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29578) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19152) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27135) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22350) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25737) * $signed(input_fmap_77[7:0]) +
	( 8'sd 118) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2540) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11523) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19844) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16055) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26957) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30544) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7997) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31251) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3660) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15663) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15139) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_95[7:0]) +
	( 10'sd 459) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31756) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9056) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17859) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16454) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11481) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7396) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28055) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3409) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27190) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10755) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14105) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2458) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7690) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9482) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14936) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5754) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13692) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8667) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21084) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26162) * $signed(input_fmap_127[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 16'd29656;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 14'd7773;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 13'd3702;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 11'd861;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 14'd6607;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 14'd8152;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 14'd4512;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 14'd7685;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 14'd5362;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 16'd22838;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 15'd16310;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 12'd1336;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 14'd4323;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 14'd6626;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 15'd14956;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 16'd24444;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 14'd7734;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 15'd11913;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 14'd6694;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 16'd27792;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 16'd17089;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 16'd27366;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 16'd23289;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 16'd22468;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 13'd2792;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 16'd26128;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 15'd8704;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 15'd12317;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 15'd13577;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 15'd13326;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 15'd14329;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 11'd1023;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 16'd28759;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 16'd18365;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 12'd1209;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 14'd5990;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 15'd15096;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 15'd11361;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 15'd10249;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 16'd25929;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 16'd25860;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 16'd26460;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 16'd16631;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 16'd23254;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 14'd7841;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 16'd24832;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 15'd15376;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 16'd24176;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 16'd27767;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 12'd1270;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 14'd7119;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 16'd19199;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 15'd9170;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 15'd10363;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 16'd20250;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 16'd19144;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 16'd16707;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 16'd20052;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 16'd24938;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 16'd18519;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 16'd16874;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 16'd20746;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 14'd7767;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 16'd23172;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 16'd21497;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 14'd6826;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 16'd32091;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 16'd30584;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 16'd29296;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 14'd4197;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 14'd8152;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 16'd22856;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 12'd1548;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 14'd6725;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 16'd25495;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 15'd12806;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 15'd15529;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 16'd28156;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 14'd4349;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 16'd23537;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 15'd13566;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 14'd5473;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 15'd13589;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 14'd4531;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 16'd22600;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 16'd31968;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 15'd14628;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 16'd32122;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 16'd26932;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 16'd26628;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 15'd11318;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 16'd29237;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 16'd21326;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 16'd25661;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 16'd20657;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 16'd18226;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 16'd28161;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 16'd30191;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 16'd26427;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 16'd31553;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 12'd1308;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 16'd28911;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 14'd5753;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 16'd21643;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 16'd21175;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 16'd27312;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 13'd3944;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 16'd18114;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 16'd23564;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 16'd18395;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 12'd1475;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 16'd17359;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 14'd4731;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 14'd6321;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 14'd4338;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 16'd18793;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 16'd17688;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 14'd5774;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 15'd10095;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 16'd24674;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 15'd9510;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 16'd21045;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 16'd25241;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 16'd28979;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 14'd4866;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 15'd9968;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 14'd4912;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 16'd26102;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[21:15]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[21:15]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[21:15]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[21:15]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[21:15]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[21:15]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[21:15]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[21:15]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[21:15]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[21:15]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[21:15]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[21:15]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[21:15]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[21:15]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[21:15]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[21:15]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[21:15]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[21:15]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[21:15]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[21:15]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[21:15]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[21:15]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[21:15]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[21:15]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[21:15]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[21:15]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[21:15]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[21:15]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[21:15]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[21:15]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[21:15]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[21:15]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[21:15]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[21:15]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[21:15]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[21:15]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[21:15]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[21:15]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[21:15]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[21:15]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[21:15]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[21:15]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[21:15]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[21:15]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[21:15]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[21:15]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[21:15]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[21:15]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[21:15]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[21:15]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[21:15]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[21:15]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[21:15]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[21:15]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[21:15]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[21:15]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[21:15]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[21:15]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[21:15]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[21:15]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[21:15]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[21:15]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[21:15]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[21:15]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[21:15]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[21:15]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[21:15]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[21:15]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[21:15]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[21:15]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[21:15]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[21:15]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[21:15]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[21:15]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[21:15]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[21:15]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[21:15]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[21:15]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[21:15]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[21:15]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[21:15]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[21:15]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[21:15]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[21:15]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[21:15]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[21:15]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[21:15]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[21:15]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[21:15]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[21:15]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[21:15]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[21:15]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[21:15]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[21:15]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[21:15]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[21:15]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[21:15]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[21:15]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[21:15]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[21:15]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[21:15]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[21:15]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[21:15]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[21:15]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[21:15]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[21:15]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[21:15]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[21:15]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[21:15]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[21:15]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[21:15]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[21:15]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[21:15]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[21:15]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[21:15]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[21:15]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[21:15]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[21:15]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[21:15]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[21:15]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[21:15]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[21:15]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[21:15]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[21:15]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[21:15]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[21:15]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[21:15]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[21:15]}} :'d6) : '0;

assign output_act = {
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
