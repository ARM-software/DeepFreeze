module conv13_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [1024-1:0] input_act,
    output logic [2048-1:0] output_act,
    output logic ready
);

logic [1024-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 16'sd 25571) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5786) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8355) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28788) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9621) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19251) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13748) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24945) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14581) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20128) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23199) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29060) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32405) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12337) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31678) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1593) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11340) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9534) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22945) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1216) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1202) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21159) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16448) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11180) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23526) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27500) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26189) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26603) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11997) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29770) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9987) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7618) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8703) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16872) * $signed(input_fmap_54[7:0]) +
	( 10'sd 274) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25224) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22836) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14208) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12101) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9044) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1076) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19703) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6029) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11670) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10203) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6109) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3952) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6893) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25788) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27037) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28234) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20383) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25431) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15831) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32664) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12610) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9290) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21669) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25663) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11807) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24164) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8691) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18871) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20180) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15401) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17847) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9306) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9950) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18741) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22903) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26671) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32197) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5995) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1859) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2268) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_123[7:0]) +
	( 10'sd 383) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10699) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25627) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24558) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 16'sd 18171) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5845) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31505) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1956) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26285) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29931) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24131) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29613) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4721) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12532) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2904) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15930) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10039) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32724) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12279) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16662) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3878) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9041) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21978) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10890) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10848) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3101) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11711) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16212) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26304) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20458) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31321) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20520) * $signed(input_fmap_49[7:0]) +
	( 8'sd 105) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2950) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6158) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23882) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8738) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1984) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32425) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18610) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6087) * $signed(input_fmap_64[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3059) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24105) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17485) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4132) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4771) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10258) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29929) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24524) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14655) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8347) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22352) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11070) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27726) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12265) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16022) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20458) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13315) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16024) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16511) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13866) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32021) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6106) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28373) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30278) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2815) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23061) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5634) * $signed(input_fmap_103[7:0]) +
	( 14'sd 8092) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31772) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4258) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3890) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3585) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12782) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20012) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10754) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4346) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31783) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11516) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2145) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_124[7:0]) +
	( 12'sd 2002) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 16'sd 22241) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8417) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32542) * $signed(input_fmap_2[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30907) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24192) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19217) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27264) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1283) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17165) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17884) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29779) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2689) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7167) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10310) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8431) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25260) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9701) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24870) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5118) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15490) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2183) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1483) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3084) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24190) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27370) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18954) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28346) * $signed(input_fmap_37[7:0]) +
	( 10'sd 417) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27959) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19357) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24893) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31684) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2891) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18841) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23915) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6895) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31020) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17077) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18344) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9260) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22982) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9499) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6888) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21291) * $signed(input_fmap_69[7:0]) +
	( 12'sd 2005) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5057) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20361) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5168) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28217) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20264) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26616) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4167) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14491) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29285) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15382) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14037) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28724) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17082) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25526) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15437) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1352) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1352) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7931) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19294) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32328) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21082) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9155) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3648) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22841) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27665) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19592) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_107[7:0]) +
	( 11'sd 850) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32145) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25604) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21657) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10311) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4833) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30610) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21904) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6439) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12339) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8244) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8013) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 16'sd 21114) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14143) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_4[7:0]) +
	( 11'sd 608) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3459) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3523) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8915) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15493) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4324) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21867) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7611) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26228) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18246) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22428) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9280) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9019) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17505) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12490) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17656) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21049) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2765) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11490) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23336) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3829) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22867) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21542) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9821) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22579) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25685) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7776) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19560) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5098) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5203) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29126) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6476) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2989) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6703) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3505) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17186) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2503) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2253) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17581) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22435) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6751) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18925) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_75[7:0]) +
	( 10'sd 446) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31435) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25092) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24545) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14614) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17713) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2591) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13561) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7513) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25379) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2698) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7667) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7810) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19202) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9260) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22841) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1867) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7185) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8348) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22466) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28742) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20601) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30408) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23009) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29851) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21324) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9991) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14809) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16003) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8275) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22874) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13695) * $signed(input_fmap_123[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27696) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29980) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 16'sd 16749) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12577) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4325) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13158) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11762) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20923) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19998) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7159) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21695) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10612) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31771) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10645) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6394) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1377) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21439) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27440) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27723) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32613) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8484) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4615) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16823) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31306) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2361) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29245) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15961) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24292) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8511) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27677) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4111) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23711) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28936) * $signed(input_fmap_43[7:0]) +
	( 9'sd 169) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12596) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25949) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31498) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8742) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17629) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13998) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1285) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1197) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17323) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18357) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25306) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9074) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7602) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_65[7:0]) +
	( 10'sd 505) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7048) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19512) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26950) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14502) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26019) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31362) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11133) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18084) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32516) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14938) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14254) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_85[7:0]) +
	( 11'sd 912) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29993) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8915) * $signed(input_fmap_89[7:0]) +
	( 10'sd 469) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28541) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32416) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7277) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21392) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10116) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29678) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23102) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32032) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25696) * $signed(input_fmap_101[7:0]) +
	( 11'sd 654) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7495) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7750) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11652) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30765) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12590) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28291) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25513) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8551) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17592) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29334) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27665) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27690) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21347) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30380) * $signed(input_fmap_121[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32749) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21331) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 15'sd 13520) * $signed(input_fmap_0[7:0]) +
	( 11'sd 840) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3996) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5950) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9580) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9598) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31843) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23824) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5266) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13198) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31428) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23806) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17587) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18734) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12137) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31967) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8316) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26922) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31148) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14025) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10286) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2194) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27471) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17573) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4949) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6343) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30716) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2352) * $signed(input_fmap_40[7:0]) +
	( 8'sd 66) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31138) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1292) * $signed(input_fmap_48[7:0]) +
	( 11'sd 514) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15508) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5111) * $signed(input_fmap_51[7:0]) +
	( 9'sd 147) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12669) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13146) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14256) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21455) * $signed(input_fmap_57[7:0]) +
	( 14'sd 8012) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13206) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16486) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12508) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28033) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1065) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9042) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10796) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29305) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31469) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_73[7:0]) +
	( 11'sd 797) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31989) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_76[7:0]) +
	( 11'sd 650) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31942) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3345) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24377) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30950) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14582) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8475) * $signed(input_fmap_92[7:0]) +
	( 11'sd 762) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5951) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25461) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28327) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28290) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18954) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31406) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31827) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25885) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30112) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3575) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25932) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8895) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16884) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15914) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31974) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 16'sd 28055) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15866) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15576) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32059) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20675) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20581) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3640) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6723) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15606) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19856) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31381) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4996) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8809) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11851) * $signed(input_fmap_20[7:0]) +
	( 6'sd 20) * $signed(input_fmap_21[7:0]) +
	( 12'sd 2035) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11648) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20153) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23113) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22493) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26699) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9015) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26486) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15357) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2925) * $signed(input_fmap_37[7:0]) +
	( 11'sd 874) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3823) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20397) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26311) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20754) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26280) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17327) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26199) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16380) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11186) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20260) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6343) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9791) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19512) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27436) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7579) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6641) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24807) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21657) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20069) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30995) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1337) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7536) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16100) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22330) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26764) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25710) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7584) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1418) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22138) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9211) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24600) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10129) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21045) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12722) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6903) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8197) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20691) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32306) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7909) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23237) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4482) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30694) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_105[7:0]) +
	( 10'sd 440) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26824) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29831) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29738) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_111[7:0]) +
	( 11'sd 906) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20829) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22988) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23207) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10161) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4675) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4118) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7362) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17219) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31153) * $signed(input_fmap_124[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5561) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 14'sd 5725) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26892) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13848) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27121) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25113) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17906) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29929) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9041) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19197) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5774) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11619) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28542) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9583) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30140) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21390) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14580) * $signed(input_fmap_27[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15571) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32152) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11523) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31372) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6957) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14984) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19710) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8957) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18181) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23697) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8488) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32060) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22084) * $signed(input_fmap_51[7:0]) +
	( 11'sd 732) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7093) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11826) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8313) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5352) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30328) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24397) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25918) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14283) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25314) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9756) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16935) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27992) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26752) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8978) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15161) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22640) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21533) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7673) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8603) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20031) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24773) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20185) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16867) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3542) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4480) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14648) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11399) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16791) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29450) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18194) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31420) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2408) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21572) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10114) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17696) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1278) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12317) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1827) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6291) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10366) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16577) * $signed(input_fmap_119[7:0]) +
	( 12'sd 2008) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20909) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6861) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 16'sd 19205) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_1[7:0]) +
	( 9'sd 233) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3288) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19728) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4243) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29330) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13890) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26940) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31954) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31035) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24512) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9572) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29888) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11487) * $signed(input_fmap_19[7:0]) +
	( 11'sd 571) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24813) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25522) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16151) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3557) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21735) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32229) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18527) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20658) * $signed(input_fmap_33[7:0]) +
	( 10'sd 385) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21960) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21765) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4711) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12291) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7660) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19066) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25760) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12825) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32020) * $signed(input_fmap_48[7:0]) +
	( 11'sd 690) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14351) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31283) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31577) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3119) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11912) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13162) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3308) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3845) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2673) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21532) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5682) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25397) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19996) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21274) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4675) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21762) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1875) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29695) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31595) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8484) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8265) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22575) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13273) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19323) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29492) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17953) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16207) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27251) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_90[7:0]) +
	( 10'sd 288) * $signed(input_fmap_91[7:0]) +
	( 11'sd 556) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3009) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15748) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1081) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2894) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2328) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26561) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7684) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15622) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14484) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3506) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27171) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8918) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28585) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_114[7:0]) +
	( 10'sd 323) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14030) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27836) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31956) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3444) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4495) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11434) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22653) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19895) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 15'sd 8518) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7067) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18865) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21402) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23287) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14610) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14284) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25031) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12964) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3826) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31211) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5918) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32709) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16717) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7984) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24560) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5651) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21802) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5058) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18200) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20926) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12344) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3970) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18109) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26343) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1872) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27196) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11016) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26335) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8582) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14838) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3258) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11218) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29144) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9511) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2496) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23519) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31419) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10234) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28704) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1871) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25730) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22136) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31323) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4478) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18949) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5832) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22009) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5382) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22562) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20065) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10388) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13577) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18053) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22789) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4821) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1917) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10518) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27371) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25702) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2249) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26568) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6913) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16484) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25070) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15151) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13381) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 16'sd 18910) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20228) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29745) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24628) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15828) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9605) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8278) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18109) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5188) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3074) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22349) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7259) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15754) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12235) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16024) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28354) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1437) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18328) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29360) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14789) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29499) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24667) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32424) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31171) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29698) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5226) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1845) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9991) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7981) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7351) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20573) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7279) * $signed(input_fmap_44[7:0]) +
	( 14'sd 8119) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29345) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23894) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23649) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17290) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17956) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5268) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11732) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16077) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21209) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26583) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_65[7:0]) +
	( 11'sd 655) * $signed(input_fmap_66[7:0]) +
	( 8'sd 83) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10521) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20216) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8130) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1465) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16884) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27211) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9511) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19001) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6847) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26918) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2409) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4270) * $signed(input_fmap_87[7:0]) +
	( 13'sd 4091) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9897) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18090) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24121) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5619) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4800) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16809) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25292) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2269) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9326) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11498) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32558) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4820) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28742) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19984) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8751) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4554) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9437) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2606) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24462) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30548) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4759) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 16'sd 16866) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_1[7:0]) +
	( 11'sd 746) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26868) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32147) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7776) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28387) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16844) * $signed(input_fmap_8[7:0]) +
	( 11'sd 726) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6241) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8407) * $signed(input_fmap_12[7:0]) +
	( 8'sd 66) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3875) * $signed(input_fmap_14[7:0]) +
	( 11'sd 969) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23551) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8664) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20590) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2519) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6636) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31582) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13787) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17586) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18123) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_25[7:0]) +
	( 11'sd 736) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1544) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28864) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1061) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25583) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23410) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10318) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28524) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11343) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16945) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26350) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5787) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11843) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26331) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5499) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5426) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6727) * $signed(input_fmap_57[7:0]) +
	( 7'sd 41) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21027) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16095) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14620) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26211) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30093) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27878) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16817) * $signed(input_fmap_74[7:0]) +
	( 11'sd 701) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27767) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21920) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5424) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21309) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14521) * $signed(input_fmap_84[7:0]) +
	( 8'sd 125) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_86[7:0]) +
	( 11'sd 544) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13614) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17359) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12309) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7889) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29465) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1482) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9968) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21864) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10337) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10169) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29570) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30457) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22389) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12972) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28712) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32635) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12459) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24822) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3463) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31014) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31240) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30474) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15816) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1205) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9281) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19619) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6591) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 16'sd 21037) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24478) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2779) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_5[7:0]) +
	( 11'sd 634) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12194) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12769) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5703) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28493) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18259) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12562) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8355) * $signed(input_fmap_18[7:0]) +
	( 11'sd 622) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23669) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9297) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14311) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4534) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23281) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9043) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1580) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23697) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19958) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5537) * $signed(input_fmap_31[7:0]) +
	( 14'sd 8151) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20927) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4497) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16038) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18308) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14586) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32049) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6992) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3958) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4609) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27749) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24008) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8502) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17354) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1549) * $signed(input_fmap_48[7:0]) +
	( 9'sd 217) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6650) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14349) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19504) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4519) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21974) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13777) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31132) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28842) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22582) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21541) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17882) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22561) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29054) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5006) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13358) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23331) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11601) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28003) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19365) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21051) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18378) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14540) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16490) * $signed(input_fmap_80[7:0]) +
	( 11'sd 764) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12030) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8466) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8789) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28867) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8199) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25875) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17280) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26972) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_95[7:0]) +
	( 10'sd 283) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6189) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_102[7:0]) +
	( 7'sd 33) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1608) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27084) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18521) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12577) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17881) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32403) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13124) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32534) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28674) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_119[7:0]) +
	( 10'sd 314) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8151) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26106) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30808) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30115) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22842) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14562) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 15'sd 12746) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4330) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19985) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32229) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16891) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32177) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26684) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23726) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27990) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13337) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16017) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9400) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7903) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3610) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15145) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14313) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30288) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27947) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6512) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7108) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21087) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31526) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4118) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9809) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21169) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15786) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4885) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5752) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22335) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4561) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7337) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2771) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31448) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30967) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21715) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27873) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26359) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9066) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21517) * $signed(input_fmap_59[7:0]) +
	( 9'sd 194) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10743) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24183) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25219) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21072) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30780) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13936) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18902) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26770) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16383) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6441) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22942) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13324) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1547) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_84[7:0]) +
	( 9'sd 234) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16843) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30731) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29048) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10090) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18612) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9706) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15079) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16417) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18582) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27182) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7653) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13438) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6333) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14259) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1316) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23878) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18298) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16923) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12868) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19454) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_118[7:0]) +
	( 9'sd 254) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2661) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10084) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10117) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30257) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12730) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 16'sd 25142) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4545) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23038) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22811) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_5[7:0]) +
	( 11'sd 908) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14698) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27325) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29257) * $signed(input_fmap_9[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15430) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22730) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27259) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30231) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20896) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9983) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30649) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10608) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4433) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2277) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10106) * $signed(input_fmap_28[7:0]) +
	( 11'sd 903) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16366) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27975) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18058) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25244) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11939) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19643) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22485) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30556) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24155) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15966) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17557) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23794) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31777) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29331) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24375) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1866) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8856) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28457) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11277) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23340) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2837) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21191) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13683) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30376) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14248) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16806) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29404) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29574) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8474) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29631) * $signed(input_fmap_82[7:0]) +
	( 9'sd 162) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23450) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2714) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23693) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22075) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24139) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1480) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19368) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24542) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26382) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29541) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16111) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3068) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26879) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7792) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17156) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10436) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11087) * $signed(input_fmap_116[7:0]) +
	( 8'sd 64) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31855) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10374) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29851) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23241) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17772) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15639) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11131) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 16'sd 18085) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12984) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16388) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18049) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31179) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16534) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22647) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5421) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2168) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5144) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9937) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4737) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15660) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5797) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6407) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25339) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13113) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15823) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13268) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18674) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32437) * $signed(input_fmap_35[7:0]) +
	( 10'sd 481) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20914) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29397) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21227) * $signed(input_fmap_41[7:0]) +
	( 10'sd 427) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21810) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13241) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9262) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18005) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7944) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19432) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10407) * $signed(input_fmap_49[7:0]) +
	( 11'sd 980) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12560) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26032) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19983) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17804) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32247) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7752) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6575) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7414) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24375) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1937) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25931) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31884) * $signed(input_fmap_67[7:0]) +
	( 11'sd 716) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22114) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22395) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13202) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31471) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29581) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8712) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16528) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1261) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20157) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26102) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1197) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23552) * $signed(input_fmap_91[7:0]) +
	( 11'sd 539) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23345) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7446) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2807) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4711) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21290) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20422) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29437) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31286) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32034) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25193) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8035) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32070) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16955) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26977) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5378) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8610) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5844) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7202) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4484) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6856) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 12'sd 1062) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20432) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32707) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21734) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6386) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13410) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18400) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30286) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16290) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17001) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5545) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_26[7:0]) +
	( 11'sd 586) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14686) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24592) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22392) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32030) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17351) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14843) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17375) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25909) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12525) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3944) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3964) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7417) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10755) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21417) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14156) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18841) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14879) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27093) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14171) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1995) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24450) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_62[7:0]) +
	( 9'sd 232) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21366) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8955) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31408) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2736) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4857) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22072) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24240) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25047) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11405) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6411) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4418) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14154) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29331) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20236) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6355) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28577) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22396) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8877) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20730) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_97[7:0]) +
	( 13'sd 4039) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29497) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23344) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23961) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22045) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8593) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8649) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20663) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18835) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8928) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12793) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3958) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25917) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30336) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8357) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15044) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16597) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2685) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 16'sd 24838) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28677) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12116) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17690) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5473) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6841) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32091) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28443) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13970) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31186) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7364) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3782) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24558) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4800) * $signed(input_fmap_16[7:0]) +
	( 10'sd 393) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3622) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4530) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4484) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17852) * $signed(input_fmap_22[7:0]) +
	( 11'sd 822) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13598) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4397) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15067) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21846) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4650) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1440) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_31[7:0]) +
	( 11'sd 813) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8951) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14373) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17242) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26843) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12355) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26099) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14000) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9098) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3682) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31998) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23160) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9180) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9345) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28059) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27060) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11769) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17579) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12542) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13039) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8459) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3117) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5106) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10803) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2398) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17842) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16501) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24336) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14841) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18429) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25835) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12216) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23890) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15167) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_87[7:0]) +
	( 10'sd 334) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30148) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14591) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9166) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26163) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20300) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17841) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26347) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1539) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28714) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23432) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23542) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13416) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24730) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7641) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32051) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9206) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24396) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20428) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22416) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20847) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31584) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29279) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15072) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7401) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19010) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10677) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7821) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 16'sd 29474) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21657) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5579) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4510) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_5[7:0]) +
	( 14'sd 8025) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5891) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14136) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13385) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20604) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31561) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26303) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29577) * $signed(input_fmap_16[7:0]) +
	( 14'sd 8101) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11747) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11302) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3588) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27078) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4416) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20217) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1701) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31676) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21482) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10477) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17009) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13115) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12915) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5687) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32138) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20138) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2899) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10414) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8281) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12028) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1483) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3795) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25684) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28362) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24445) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3930) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21990) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6231) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29947) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9963) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22488) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2101) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18406) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16580) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29541) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27456) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30700) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31019) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_73[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29247) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22184) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8424) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18574) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14584) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5491) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20798) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20111) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24954) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21580) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4250) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1786) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11995) * $signed(input_fmap_96[7:0]) +
	( 13'sd 4072) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8649) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_102[7:0]) +
	( 11'sd 971) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13862) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10071) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9734) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28024) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18523) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28966) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16447) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3292) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2362) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20665) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27223) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29167) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18125) * $signed(input_fmap_124[7:0]) +
	( 10'sd 264) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 16'sd 30052) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2617) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13500) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27334) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15439) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27324) * $signed(input_fmap_5[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17865) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12744) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25613) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17923) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16406) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11131) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26669) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3164) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26051) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13597) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2128) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15689) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6486) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24415) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19604) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20878) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19692) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12951) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14511) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15580) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24905) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10598) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18670) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13217) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26451) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30718) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17471) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15582) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20735) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27170) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_64[7:0]) +
	( 10'sd 343) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7212) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15762) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27887) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22310) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23687) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3331) * $signed(input_fmap_77[7:0]) +
	( 12'sd 2014) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2050) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29495) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30260) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9902) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29534) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12845) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_89[7:0]) +
	( 11'sd 863) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26665) * $signed(input_fmap_91[7:0]) +
	( 13'sd 4039) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17892) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26846) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9662) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29584) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13516) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30168) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21927) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9443) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20688) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16818) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28337) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31001) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3729) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16248) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_112[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16588) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8662) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22861) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32230) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2920) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20949) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6729) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 16'sd 20746) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3431) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15099) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1155) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10222) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15367) * $signed(input_fmap_5[7:0]) +
	( 10'sd 466) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5709) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5634) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7638) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3034) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10464) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30162) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23877) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2433) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24826) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13193) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24388) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15552) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12782) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20128) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4655) * $signed(input_fmap_25[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_27[7:0]) +
	( 11'sd 894) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14578) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30814) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16111) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31219) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8850) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28219) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16752) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22271) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7535) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12463) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16884) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29421) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25805) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15201) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22003) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21654) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32029) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8437) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21113) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31965) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25161) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_64[7:0]) +
	( 13'sd 4016) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28858) * $signed(input_fmap_67[7:0]) +
	( 10'sd 449) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10739) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22788) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8804) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14957) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1442) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7282) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9721) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15797) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28467) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14196) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_82[7:0]) +
	( 11'sd 943) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28766) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27798) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27560) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16138) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25235) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10742) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11618) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28205) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21378) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2122) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9402) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25313) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31200) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12469) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23301) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23137) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7824) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4717) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4437) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14582) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4115) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11647) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16332) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_114[7:0]) +
	( 6'sd 16) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8540) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9234) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13966) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16589) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10828) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30271) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23511) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23917) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16149) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 16'sd 26678) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29439) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18471) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25804) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2654) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4804) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26246) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9647) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_12[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7880) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16211) * $signed(input_fmap_15[7:0]) +
	( 9'sd 153) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31162) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21538) * $signed(input_fmap_20[7:0]) +
	( 13'sd 4060) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11117) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3474) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6413) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9409) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11355) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25739) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20057) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12139) * $signed(input_fmap_41[7:0]) +
	( 10'sd 444) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1937) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26545) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2975) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23805) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26395) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14099) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_51[7:0]) +
	( 13'sd 4039) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14535) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_55[7:0]) +
	( 13'sd 4061) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2860) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19373) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25344) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9102) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15385) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6257) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29085) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22262) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10551) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5572) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5959) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1125) * $signed(input_fmap_72[7:0]) +
	( 10'sd 320) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30602) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14261) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18960) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29448) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_82[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4731) * $signed(input_fmap_84[7:0]) +
	( 11'sd 684) * $signed(input_fmap_85[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7064) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1943) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25904) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23890) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17701) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21633) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9986) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19136) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30145) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7255) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5596) * $signed(input_fmap_98[7:0]) +
	( 13'sd 4087) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3711) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25064) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31747) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2422) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4729) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_109[7:0]) +
	( 11'sd 517) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15567) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4933) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21462) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3723) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_118[7:0]) +
	( 11'sd 812) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32008) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10063) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25769) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29966) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32662) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11660) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 15'sd 10414) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29279) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31043) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19644) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14433) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5964) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31465) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12408) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29976) * $signed(input_fmap_10[7:0]) +
	( 10'sd 510) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17036) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17777) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31392) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3607) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20235) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_20[7:0]) +
	( 11'sd 912) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27480) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12805) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3983) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_27[7:0]) +
	( 11'sd 897) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2847) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5259) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14467) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29812) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25987) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13758) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10067) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12861) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6621) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_42[7:0]) +
	( 11'sd 600) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6909) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31806) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27660) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6932) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23529) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6650) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11313) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10697) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20532) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1829) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27226) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_60[7:0]) +
	( 11'sd 802) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6097) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12289) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6715) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17649) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22148) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2125) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5778) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8161) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14208) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15793) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17306) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9302) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4789) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4885) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11675) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_89[7:0]) +
	( 12'sd 2046) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29497) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19055) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24280) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6701) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17042) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32448) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10627) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16536) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5124) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3720) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13892) * $signed(input_fmap_110[7:0]) +
	( 15'sd 16341) * $signed(input_fmap_111[7:0]) +
	( 12'sd 2010) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23169) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31937) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23054) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19681) * $signed(input_fmap_120[7:0]) +
	( 9'sd 238) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6786) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6015) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21003) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31710) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 16'sd 18673) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13747) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3207) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15476) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30224) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22887) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24630) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26084) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21479) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8451) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1469) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8705) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25568) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24871) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7397) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14053) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19150) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23047) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25599) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2724) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6434) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14655) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11961) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23267) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25984) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21504) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2454) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27206) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6630) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20925) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3667) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16218) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11499) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15890) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23516) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19569) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32052) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9408) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_52[7:0]) +
	( 4'sd 5) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25719) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5289) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1857) * $signed(input_fmap_57[7:0]) +
	( 9'sd 217) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17993) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17707) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15099) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11191) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1441) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19253) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15985) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17192) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15034) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14346) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16249) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26661) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_76[7:0]) +
	( 8'sd 126) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12800) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2079) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17933) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23920) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8797) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25104) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21538) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6733) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32694) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_90[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10696) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27811) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31201) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8328) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31481) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26662) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13113) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10605) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11886) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13444) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30035) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23075) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28666) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23852) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27082) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19536) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18098) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7947) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25216) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 15'sd 8734) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27223) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9638) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11588) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30122) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3424) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11191) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28652) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23036) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8338) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28730) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_20[7:0]) +
	( 9'sd 190) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21112) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31201) * $signed(input_fmap_23[7:0]) +
	( 11'sd 812) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32697) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26714) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7541) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_32[7:0]) +
	( 10'sd 489) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30637) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11551) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23986) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29866) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21330) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6235) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29724) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14306) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1540) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1503) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26113) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24357) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8357) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27104) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10583) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1858) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21679) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22048) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21716) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_74[7:0]) +
	( 11'sd 622) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1440) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27901) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8870) * $signed(input_fmap_78[7:0]) +
	( 13'sd 4041) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18083) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26663) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24658) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32260) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10736) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17575) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10695) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2496) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29973) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24678) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22838) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15990) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20735) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3073) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23800) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30218) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7459) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23860) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17071) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22914) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28482) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_113[7:0]) +
	( 11'sd 954) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31412) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12395) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2147) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3571) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10772) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3495) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30150) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15303) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28264) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26015) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1822) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 16'sd 17657) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_1[7:0]) +
	( 11'sd 961) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26436) * $signed(input_fmap_3[7:0]) +
	( 14'sd 8101) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11455) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7843) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30422) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8023) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7422) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3074) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21631) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20272) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6932) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12062) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16972) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15499) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27395) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28304) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32097) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31497) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7345) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13762) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15871) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30277) * $signed(input_fmap_33[7:0]) +
	( 11'sd 654) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18429) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18952) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12260) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30553) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4142) * $signed(input_fmap_39[7:0]) +
	( 11'sd 592) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26029) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_42[7:0]) +
	( 10'sd 260) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25056) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32018) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12139) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9931) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11463) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9133) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29334) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7394) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2107) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14023) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5690) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11314) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9914) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30440) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5049) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11765) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7611) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17930) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20057) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6932) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19380) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6437) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26120) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26890) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11854) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17268) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19324) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17721) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1472) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9679) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10584) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29081) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21366) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14818) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24166) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17495) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23025) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24480) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23923) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18040) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20943) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14559) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4706) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23984) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26576) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2347) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25169) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15986) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21574) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22990) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32558) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 15'sd 14489) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24731) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32170) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3461) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19295) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4985) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12386) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3059) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17086) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28273) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25360) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28289) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32184) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23655) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27059) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32200) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13241) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16409) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15674) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6262) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8752) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18899) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26484) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29357) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4327) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16414) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_38[7:0]) +
	( 11'sd 562) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5192) * $signed(input_fmap_41[7:0]) +
	( 9'sd 249) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19713) * $signed(input_fmap_43[7:0]) +
	( 10'sd 425) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10235) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25709) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13828) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15850) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18068) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11330) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5879) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22371) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2117) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18050) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7315) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17417) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12034) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17164) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27696) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19568) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6579) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30511) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9904) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5351) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17406) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12491) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9924) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9034) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11714) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23324) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29604) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24680) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12408) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18441) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24306) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10210) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4374) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6179) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20046) * $signed(input_fmap_106[7:0]) +
	( 11'sd 770) * $signed(input_fmap_107[7:0]) +
	( 10'sd 488) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6395) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10514) * $signed(input_fmap_110[7:0]) +
	( 11'sd 811) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32488) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3753) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8701) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9636) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24180) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20461) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1332) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6284) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11610) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14017) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20342) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 16'sd 23974) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24888) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24411) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25478) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32646) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18942) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27686) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30190) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7615) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22328) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30003) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13789) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2436) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22870) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30617) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18338) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8354) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7041) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25493) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19585) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17567) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23596) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20260) * $signed(input_fmap_36[7:0]) +
	( 11'sd 1012) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27738) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22158) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4200) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21708) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20536) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6343) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6558) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18806) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20159) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5594) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20770) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18159) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14716) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14890) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23046) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22311) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14765) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9867) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22148) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29685) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18502) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11158) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31981) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20050) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2359) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1266) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22800) * $signed(input_fmap_90[7:0]) +
	( 13'sd 4060) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10811) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13692) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11601) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21183) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2089) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26068) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28554) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13888) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7566) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5737) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28967) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7716) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14725) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25873) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14439) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25670) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21107) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10832) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22024) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26073) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30959) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23017) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16226) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24547) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16999) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 14'sd 7485) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26063) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6076) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26470) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29805) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17222) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20675) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2337) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9470) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29418) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8765) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26763) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28410) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1048) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31626) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6373) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12719) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16932) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20764) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22541) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31291) * $signed(input_fmap_34[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9163) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7036) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32040) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17366) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20714) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8658) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26320) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8591) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14794) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17499) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27240) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20347) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15012) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8853) * $signed(input_fmap_51[7:0]) +
	( 13'sd 4021) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2925) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22537) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21187) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14324) * $signed(input_fmap_56[7:0]) +
	( 11'sd 878) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8578) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16962) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18143) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16855) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24279) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7037) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14675) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18741) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4205) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2166) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4668) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9394) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31303) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31593) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28491) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9021) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24904) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22818) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13985) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9131) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26515) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5916) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20361) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14402) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3344) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1406) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2501) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28153) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16279) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4480) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2631) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16070) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32338) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32246) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13814) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6579) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29510) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10406) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29041) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20227) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9828) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21771) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20160) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11873) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 16'sd 18971) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3128) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19119) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15352) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10334) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32664) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31974) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29234) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14144) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23359) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27555) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11937) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30873) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2160) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17763) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7324) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27622) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15255) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28559) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15985) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31106) * $signed(input_fmap_27[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28755) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21400) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31531) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19058) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11949) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23184) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10320) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23246) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31187) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14380) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28011) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12827) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19746) * $signed(input_fmap_51[7:0]) +
	( 11'sd 748) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5504) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7404) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16059) * $signed(input_fmap_55[7:0]) +
	( 6'sd 25) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20299) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5180) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31810) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4831) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1731) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13061) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4444) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28254) * $signed(input_fmap_66[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30989) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30710) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29728) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8465) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18910) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3259) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31813) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31738) * $signed(input_fmap_82[7:0]) +
	( 9'sd 194) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_84[7:0]) +
	( 8'sd 95) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2244) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24022) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28177) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12092) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5409) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17158) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_96[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16546) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_101[7:0]) +
	( 11'sd 941) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27668) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_105[7:0]) +
	( 11'sd 1022) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26497) * $signed(input_fmap_107[7:0]) +
	( 10'sd 452) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10406) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9325) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22113) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_115[7:0]) +
	( 8'sd 70) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18122) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9763) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_121[7:0]) +
	( 9'sd 180) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26509) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5048) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12650) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 16'sd 25390) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17248) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11253) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5736) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27026) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32539) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23487) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29053) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4490) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28472) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28847) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18204) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18299) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3561) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7341) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19752) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2365) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6797) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1891) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6717) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22706) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14603) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20118) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25944) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6083) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19384) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17487) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22353) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30900) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29587) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32417) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4294) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2237) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28720) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31278) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28317) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30397) * $signed(input_fmap_63[7:0]) +
	( 7'sd 62) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13646) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26573) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20533) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15214) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31926) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6136) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27232) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10462) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8250) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7583) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22415) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29834) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12947) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18647) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25187) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24299) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27947) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9612) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9104) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9086) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5545) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16075) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1584) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21293) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32049) * $signed(input_fmap_106[7:0]) +
	( 11'sd 716) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29226) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17620) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25632) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6635) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22570) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18027) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_115[7:0]) +
	( 10'sd 381) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32198) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12270) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23959) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11197) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22148) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 14'sd 5337) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9924) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7352) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11864) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32700) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12752) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23538) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4396) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16823) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19897) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24363) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2317) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31321) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28988) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30769) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31265) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21871) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20938) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14401) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29669) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6068) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26002) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11754) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25813) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7353) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30023) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11458) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31673) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2341) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26474) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12093) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_50[7:0]) +
	( 15'sd 16318) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11438) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12181) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10079) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10095) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13942) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18611) * $signed(input_fmap_58[7:0]) +
	( 11'sd 554) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9324) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4108) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26836) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27999) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6368) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23818) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14535) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22169) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22711) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2754) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22760) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5670) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24635) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27387) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28346) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24268) * $signed(input_fmap_79[7:0]) +
	( 10'sd 281) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8997) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32456) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10134) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18472) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7310) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14045) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12067) * $signed(input_fmap_93[7:0]) +
	( 11'sd 906) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17762) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31377) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24631) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5247) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18417) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_102[7:0]) +
	( 11'sd 904) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8555) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14634) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22441) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11815) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21029) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4430) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3221) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16561) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22628) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1585) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28629) * $signed(input_fmap_124[7:0]) +
	( 12'sd 2037) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24640) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 15'sd 9527) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12050) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8958) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9805) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11637) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29457) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16931) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22121) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14451) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12080) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13927) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12320) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28269) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2555) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23865) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26732) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1609) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27861) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18549) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18502) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18996) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2325) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32164) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26173) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9473) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21191) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17903) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7014) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9418) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2089) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21692) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22987) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20971) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9296) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23924) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9623) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23282) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25938) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27707) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5039) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30400) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30005) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9151) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25399) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11309) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19160) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29780) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1224) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3441) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23338) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29324) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22393) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27985) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7776) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8219) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9049) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11712) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6025) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18496) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18426) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32765) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14236) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32411) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 16'sd 20820) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12344) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17927) * $signed(input_fmap_2[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5882) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20798) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5210) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25647) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32373) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24100) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18337) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11075) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7863) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9520) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14950) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6539) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15539) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28260) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25305) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31306) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17639) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27220) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10472) * $signed(input_fmap_37[7:0]) +
	( 11'sd 556) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4363) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17973) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20471) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10170) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1125) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3100) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29966) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15408) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14894) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14114) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8892) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18948) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7405) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29228) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3587) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13915) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12769) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22462) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11536) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2544) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25621) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31569) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15336) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6632) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16858) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1633) * $signed(input_fmap_78[7:0]) +
	( 6'sd 23) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2188) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22275) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25674) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9970) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25491) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6908) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9066) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12900) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18585) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15513) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13169) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29187) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2452) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31524) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25419) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13247) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7890) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20663) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10672) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10079) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4608) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30269) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24554) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30529) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29642) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3120) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12192) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 15'sd 13217) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1542) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27418) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28994) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32479) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17595) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1358) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13204) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4920) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27094) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1098) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27437) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8971) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2455) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16804) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25540) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2582) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8535) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21502) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4689) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13693) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6327) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4517) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32587) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30385) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22636) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_38[7:0]) +
	( 11'sd 846) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24358) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11123) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25870) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24801) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15783) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18404) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_51[7:0]) +
	( 10'sd 463) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1426) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10675) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1286) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26350) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15695) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3112) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9160) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8485) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2232) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4412) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26670) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30230) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20005) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31679) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6517) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30121) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12665) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13900) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14740) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3215) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4356) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15115) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14291) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28199) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30097) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29313) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10518) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18278) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10697) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18299) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16737) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5528) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24670) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6253) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24222) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31606) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1997) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24782) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17319) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14357) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22227) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30100) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22747) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14894) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24377) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18507) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10890) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11954) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12729) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 15'sd 13706) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19022) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17891) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32550) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3663) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22848) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7832) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12331) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6560) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5103) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12326) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7253) * $signed(input_fmap_16[7:0]) +
	( 11'sd 653) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27378) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3071) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23761) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_25[7:0]) +
	( 11'sd 846) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15732) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7584) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21746) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20580) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10627) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31941) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27044) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30407) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13591) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21363) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9947) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3672) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14705) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12080) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31560) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9471) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8448) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23676) * $signed(input_fmap_55[7:0]) +
	( 13'sd 4089) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12695) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10002) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26739) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26617) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30094) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17803) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24285) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9451) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13790) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4316) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7065) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6706) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8788) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23607) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26755) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27985) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9889) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8913) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16079) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18752) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27499) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30157) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3788) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20492) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1563) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9680) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25455) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6805) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29524) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28144) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18866) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9853) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19150) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16660) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10659) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13797) * $signed(input_fmap_122[7:0]) +
	( 11'sd 556) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6465) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4860) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 16'sd 16384) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28563) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21663) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26143) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7086) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3773) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23196) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1328) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7385) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26599) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18044) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30690) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22282) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7525) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1140) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32075) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9043) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25930) * $signed(input_fmap_26[7:0]) +
	( 11'sd 656) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3746) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23162) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29237) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5968) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19206) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29652) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4446) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19736) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28159) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9136) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17694) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1384) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30277) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10140) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8676) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19903) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4429) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17318) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13745) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13985) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13895) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17465) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24072) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12535) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12547) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22903) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4422) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22261) * $signed(input_fmap_67[7:0]) +
	( 10'sd 351) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10790) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16298) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4777) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4647) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24527) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21757) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13421) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7361) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3986) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28874) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32549) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1512) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13205) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19984) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18189) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12793) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25547) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7025) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16642) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18268) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7005) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22141) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24950) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11418) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2898) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16103) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3491) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14385) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29442) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6990) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8032) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2855) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6804) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28031) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2168) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11927) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18745) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 15'sd 10541) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22354) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1843) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4475) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16146) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2577) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14776) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20474) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31252) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22501) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6683) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4696) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2389) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1984) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26272) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4563) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6993) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27938) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23517) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27166) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29280) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6450) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24001) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10135) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10936) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12932) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12375) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3934) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5489) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1030) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10964) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22475) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23356) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24725) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16567) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26059) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29433) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24651) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30474) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15328) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1930) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18241) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11726) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32324) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5963) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14956) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9985) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_65[7:0]) +
	( 10'sd 302) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30140) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29814) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17507) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_70[7:0]) +
	( 11'sd 538) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18468) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21855) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24140) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3684) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23198) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23371) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6491) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32409) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19134) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25119) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7389) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3024) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_88[7:0]) +
	( 9'sd 204) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25690) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25818) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9201) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18935) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22829) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3546) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2751) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11304) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1447) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13852) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4493) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8580) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5879) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25594) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26145) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9252) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25707) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8855) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10526) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21929) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23913) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21055) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32662) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26458) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 16'sd 18840) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22731) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18590) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26832) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_8[7:0]) +
	( 8'sd 67) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27657) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8795) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5631) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22479) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13633) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18535) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27562) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10265) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5976) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3383) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20756) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20866) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20933) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28983) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20966) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16144) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18188) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31064) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32718) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16354) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6902) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6808) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7910) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30152) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29722) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1389) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10951) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5049) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22544) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7814) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18823) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10940) * $signed(input_fmap_60[7:0]) +
	( 11'sd 551) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8209) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24746) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5670) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22042) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15098) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2956) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21013) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32589) * $signed(input_fmap_69[7:0]) +
	( 13'sd 4050) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7346) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2250) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16942) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19637) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27247) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11310) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24495) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10124) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28898) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17532) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21974) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17166) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21537) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15148) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29314) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6109) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4527) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25493) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21462) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16917) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20578) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23944) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32364) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25538) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15965) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19088) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6185) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2238) * $signed(input_fmap_117[7:0]) +
	( 11'sd 564) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13927) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7002) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1199) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9666) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8211) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 16'sd 23474) * $signed(input_fmap_0[7:0]) +
	( 11'sd 606) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23237) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9554) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11268) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_7[7:0]) +
	( 11'sd 751) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14102) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5116) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7490) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25570) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21179) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22902) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30857) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13198) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8680) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32262) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1270) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26657) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27762) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32615) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27095) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28882) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3175) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24635) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31394) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25735) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24419) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25506) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30086) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25940) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23606) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24017) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16643) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20258) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23314) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19885) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14684) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18725) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1901) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22932) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15982) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2918) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3248) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29766) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28365) * $signed(input_fmap_69[7:0]) +
	( 11'sd 678) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6873) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19742) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31543) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29442) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29639) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5896) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28654) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23350) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15906) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11071) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8332) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24401) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13567) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28244) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6061) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2144) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12281) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9569) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8959) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31070) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10891) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6614) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1024) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18711) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13587) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29334) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12552) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27127) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13548) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31531) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24788) * $signed(input_fmap_113[7:0]) +
	( 10'sd 443) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26327) * $signed(input_fmap_115[7:0]) +
	( 9'sd 186) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17558) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24084) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30125) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29427) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26651) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18529) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 15'sd 8835) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26622) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16881) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16763) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_5[7:0]) +
	( 8'sd 113) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28677) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29564) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5344) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6433) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13374) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15809) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8776) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17477) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20785) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16518) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15628) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8041) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25577) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14021) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25336) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11737) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21714) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27450) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3480) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11801) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12715) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15100) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28884) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7155) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20635) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25300) * $signed(input_fmap_55[7:0]) +
	( 11'sd 844) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9456) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17712) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5153) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11598) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20422) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12860) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18055) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12948) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23174) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4930) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23856) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22872) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14403) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15271) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6070) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10357) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15388) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13987) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10519) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13862) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8715) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18116) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13859) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9439) * $signed(input_fmap_89[7:0]) +
	( 11'sd 594) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25342) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28888) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24410) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28635) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30993) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3254) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17566) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7479) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8208) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20524) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17050) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5219) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21770) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22669) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22183) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16565) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6106) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32396) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5497) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30566) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13753) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23729) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3680) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20901) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 15'sd 15829) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7650) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13040) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26446) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17931) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20014) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23031) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9756) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29204) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14564) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18947) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16966) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20997) * $signed(input_fmap_20[7:0]) +
	( 11'sd 852) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19981) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28349) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8510) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10948) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30833) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11396) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30082) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24084) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13564) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8346) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19252) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7759) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2596) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20953) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17701) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21727) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14033) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10948) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5364) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26262) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17433) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3381) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32583) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31922) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16806) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13625) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32497) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2171) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12535) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27869) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3743) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5865) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19557) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13374) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27701) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16232) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10438) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26193) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27028) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5142) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25647) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3251) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5381) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29072) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1289) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13593) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25276) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18075) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1402) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1902) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20927) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_97[7:0]) +
	( 10'sd 358) * $signed(input_fmap_98[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_100[7:0]) +
	( 11'sd 688) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14882) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3917) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20685) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15883) * $signed(input_fmap_108[7:0]) +
	( 13'sd 4056) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16061) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3458) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7267) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27068) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20459) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6210) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13062) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32523) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30548) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15016) * $signed(input_fmap_125[7:0]) +
	( 6'sd 21) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 15'sd 13420) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15344) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7481) * $signed(input_fmap_3[7:0]) +
	( 10'sd 327) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20922) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19632) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27573) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32371) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21032) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21518) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14376) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9381) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15612) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27916) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25711) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11167) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18664) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15970) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6560) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29885) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7928) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11307) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9299) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16273) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10333) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25606) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20620) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12157) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11156) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21578) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9096) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32652) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24570) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5593) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23082) * $signed(input_fmap_51[7:0]) +
	( 11'sd 879) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10862) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7557) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27550) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21700) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23395) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26865) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21335) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6085) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10937) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25549) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7680) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29942) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31604) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29096) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20072) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24037) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6441) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24928) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_79[7:0]) +
	( 10'sd 505) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24216) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3250) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32157) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24960) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12032) * $signed(input_fmap_87[7:0]) +
	( 8'sd 82) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16739) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14968) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17870) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6478) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16270) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22892) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11326) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28460) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26278) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_107[7:0]) +
	( 11'sd 793) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22929) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15863) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28804) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14192) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6622) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20500) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6400) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8852) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18286) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14101) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_123[7:0]) +
	( 12'sd 2002) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19910) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 14'sd 6531) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30787) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21370) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3226) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9782) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12429) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4865) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6691) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16556) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24777) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10629) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_13[7:0]) +
	( 7'sd 57) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22915) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8581) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18790) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15564) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21584) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22886) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6189) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13515) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2292) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14521) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10742) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30860) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25024) * $signed(input_fmap_37[7:0]) +
	( 11'sd 909) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18932) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5364) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3607) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22959) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11157) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5253) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3656) * $signed(input_fmap_47[7:0]) +
	( 13'sd 4078) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28361) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16554) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17995) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2983) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11874) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11078) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7914) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29551) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28173) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16060) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3346) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10297) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20178) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6246) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7781) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25940) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8306) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32183) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8301) * $signed(input_fmap_77[7:0]) +
	( 8'sd 84) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5223) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20232) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_82[7:0]) +
	( 10'sd 420) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14838) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20783) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10733) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22799) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20423) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14284) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28987) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1421) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23059) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14972) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22560) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22361) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20744) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15365) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22649) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15875) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23615) * $signed(input_fmap_106[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11752) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19910) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1071) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18942) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21738) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15606) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14603) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24452) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7420) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15085) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29249) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20583) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3175) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 14'sd 4748) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10518) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15248) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7572) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15009) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24573) * $signed(input_fmap_9[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22176) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16019) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2539) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3502) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18541) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19872) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14998) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11443) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10023) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31908) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_25[7:0]) +
	( 8'sd 69) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22749) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25227) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2830) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19899) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19802) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5692) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25876) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8323) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26557) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16312) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8538) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29309) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13550) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2252) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10076) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24779) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10823) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32115) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21229) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11489) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13981) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12440) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32707) * $signed(input_fmap_64[7:0]) +
	( 6'sd 23) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32705) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5634) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16657) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1821) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3871) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17063) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24785) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32407) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21469) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29778) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7691) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31506) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17276) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3424) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32019) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5682) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27973) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31285) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18772) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17074) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2923) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27024) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12959) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16963) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24698) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15747) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26603) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21884) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14644) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16390) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6406) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27265) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1169) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20141) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15032) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3310) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26015) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23464) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7889) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13666) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27190) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32662) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 16'sd 28823) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29698) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17861) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18744) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1998) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28786) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29728) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9088) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6853) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32439) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19383) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19938) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8892) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27526) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32407) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9418) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16232) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7757) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15301) * $signed(input_fmap_24[7:0]) +
	( 7'sd 41) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21165) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1370) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29764) * $signed(input_fmap_33[7:0]) +
	( 10'sd 467) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15226) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29828) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9017) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23960) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2074) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23649) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25137) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27985) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7878) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19837) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28563) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19460) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32070) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3908) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30513) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20231) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4723) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19611) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29894) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29763) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18039) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2819) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18767) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29175) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27806) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16253) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27278) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10582) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11975) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30700) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1833) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22081) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23598) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31824) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23599) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12000) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2459) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19402) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2314) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11239) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24687) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28018) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25774) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10969) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12220) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30189) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12043) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27068) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20303) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9660) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20309) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22347) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12015) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18717) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27958) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16233) * $signed(input_fmap_117[7:0]) +
	( 13'sd 4053) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23476) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21215) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22574) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22771) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 16'sd 22117) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2171) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30738) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22799) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5907) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13920) * $signed(input_fmap_7[7:0]) +
	( 13'sd 4050) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22497) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1319) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29042) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5800) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14596) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9413) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28785) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19458) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29896) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10255) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12160) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18899) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5141) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_25[7:0]) +
	( 11'sd 583) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23657) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5302) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12339) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31263) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25540) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17044) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29093) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18794) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16087) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22803) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20753) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19505) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17984) * $signed(input_fmap_44[7:0]) +
	( 11'sd 773) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9894) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12402) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21457) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3414) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5519) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18079) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7318) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22611) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5702) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13617) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14281) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32055) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31873) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27616) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15125) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31912) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31203) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21865) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24662) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17518) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20354) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11365) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25022) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1370) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28799) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4783) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20396) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25477) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30825) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21950) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32490) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15697) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1753) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17888) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18822) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18006) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_102[7:0]) +
	( 8'sd 122) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17603) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14501) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11269) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15219) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9622) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12739) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25726) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30771) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32706) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29831) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7427) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2827) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30221) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4413) * $signed(input_fmap_124[7:0]) +
	( 10'sd 395) * $signed(input_fmap_125[7:0]) +
	( 14'sd 8164) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17735) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 14'sd 4557) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9783) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19017) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21501) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12975) * $signed(input_fmap_7[7:0]) +
	( 8'sd 77) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5554) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22119) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19775) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22398) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23576) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24793) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31655) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14191) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23173) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15247) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3313) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18844) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18252) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11425) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27747) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4186) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21708) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22511) * $signed(input_fmap_48[7:0]) +
	( 11'sd 972) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22065) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13415) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20339) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8763) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31572) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7464) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9546) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11990) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16697) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25963) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5339) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22460) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2152) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10736) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30726) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15047) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13768) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28439) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10620) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14989) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5846) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31445) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7283) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3878) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10636) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31510) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14781) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16284) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14811) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16162) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14045) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3691) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4682) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6951) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15546) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10397) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8776) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19649) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26481) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30119) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14883) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10808) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23273) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32380) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5036) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4935) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4845) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8720) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29907) * $signed(input_fmap_120[7:0]) +
	( 11'sd 992) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25832) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17282) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13360) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 16'sd 23763) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15931) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26879) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27343) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32301) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6670) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18898) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19903) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11753) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20625) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12323) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22098) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3263) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3225) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7594) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18534) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17804) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2235) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26265) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20721) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5224) * $signed(input_fmap_46[7:0]) +
	( 11'sd 639) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6180) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19121) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2453) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14893) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27176) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12934) * $signed(input_fmap_55[7:0]) +
	( 10'sd 394) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28229) * $signed(input_fmap_57[7:0]) +
	( 9'sd 144) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30857) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14470) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26931) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1264) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6150) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17945) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27463) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10684) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9769) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19391) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20656) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31990) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32353) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30122) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31545) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9668) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14413) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6222) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29030) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29067) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2523) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27789) * $signed(input_fmap_89[7:0]) +
	( 11'sd 916) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11974) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22524) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16990) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31600) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31237) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_103[7:0]) +
	( 11'sd 740) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14642) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12257) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2371) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13652) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23264) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8634) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18057) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7476) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24407) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24663) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19934) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4612) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11185) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15541) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 13'sd 2612) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29067) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31443) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15741) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12990) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13275) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10153) * $signed(input_fmap_8[7:0]) +
	( 10'sd 348) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10484) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12478) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12980) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26792) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5589) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23213) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20009) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16006) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18219) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16160) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2148) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23610) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10894) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25121) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32230) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28616) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5481) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20761) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3030) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21842) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10998) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19909) * $signed(input_fmap_44[7:0]) +
	( 10'sd 463) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10276) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30876) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5450) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7041) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3722) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30431) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19548) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31152) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7320) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15965) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20603) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24808) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2988) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5832) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11189) * $signed(input_fmap_68[7:0]) +
	( 11'sd 861) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31421) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5273) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26989) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18517) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2816) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26502) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9367) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22537) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13090) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31023) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19798) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1205) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11466) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3009) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4172) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27346) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1083) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7179) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9872) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3026) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29443) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17910) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26669) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17196) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7537) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19174) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23052) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16290) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11424) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26295) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31136) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20984) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27206) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23248) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10329) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25158) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27593) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27242) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3822) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 15'sd 11283) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19701) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29444) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16798) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32027) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27909) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25434) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25903) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15460) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19573) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6077) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12630) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27729) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5536) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32429) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14094) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28283) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8750) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30814) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10010) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15683) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8783) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13411) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5031) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31364) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7309) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16956) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15692) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27107) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_46[7:0]) +
	( 13'sd 4061) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16802) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_49[7:0]) +
	( 11'sd 528) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28248) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24775) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21166) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8716) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29539) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27315) * $signed(input_fmap_61[7:0]) +
	( 9'sd 152) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21757) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23847) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12627) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9209) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28588) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_73[7:0]) +
	( 4'sd 5) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2710) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21139) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2345) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1082) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17532) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21406) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22859) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29503) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4418) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5868) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1550) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13285) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6613) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_92[7:0]) +
	( 11'sd 972) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27060) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4790) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7914) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26821) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28314) * $signed(input_fmap_99[7:0]) +
	( 12'sd 2002) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5677) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9867) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15403) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19841) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30384) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6430) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10130) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21854) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18904) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20433) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32004) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23817) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4874) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1788) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28776) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 15'sd 14095) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17670) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31586) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19469) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23530) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32070) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10714) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18055) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1632) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4752) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7166) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24625) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6372) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15096) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21280) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16921) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21880) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9928) * $signed(input_fmap_18[7:0]) +
	( 11'sd 903) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30012) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_23[7:0]) +
	( 11'sd 670) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2168) * $signed(input_fmap_25[7:0]) +
	( 10'sd 427) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3231) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8306) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11774) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25463) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12331) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6896) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14193) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5994) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4181) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3526) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21927) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23572) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22679) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28122) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7431) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27467) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17542) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20979) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19558) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24937) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13182) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20630) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7666) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3836) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25261) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24070) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29893) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15881) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4825) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16190) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16986) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2427) * $signed(input_fmap_76[7:0]) +
	( 11'sd 530) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15927) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3328) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12496) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28492) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13889) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23116) * $signed(input_fmap_88[7:0]) +
	( 10'sd 383) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32296) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4778) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_93[7:0]) +
	( 11'sd 520) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24698) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26014) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25410) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7851) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29121) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10310) * $signed(input_fmap_103[7:0]) +
	( 11'sd 692) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20862) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11945) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32488) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20162) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26206) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9773) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9539) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10485) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4318) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13352) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2680) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16297) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10579) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 13'sd 2141) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11495) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13837) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13354) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25757) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30462) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14021) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10744) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31789) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32764) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27170) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20896) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21220) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10569) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31884) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19466) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28278) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11834) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8409) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31398) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6806) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20574) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30224) * $signed(input_fmap_34[7:0]) +
	( 9'sd 197) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5474) * $signed(input_fmap_36[7:0]) +
	( 11'sd 863) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11815) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31861) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20521) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26059) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15805) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16847) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15676) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24091) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4169) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28364) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24859) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28958) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31367) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1281) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19935) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25844) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7339) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11730) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27387) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9058) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12254) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26348) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6990) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_77[7:0]) +
	( 13'sd 4037) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20659) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11125) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23069) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6805) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26801) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29595) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29652) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26587) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18784) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25345) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21383) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2667) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20176) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15421) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20389) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3345) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13047) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4402) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30411) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26113) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12538) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7073) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16996) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22819) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29213) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14948) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 16'sd 29332) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8777) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9024) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32687) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8557) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_6[7:0]) +
	( 11'sd 639) * $signed(input_fmap_7[7:0]) +
	( 11'sd 984) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12595) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12790) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25083) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4574) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3988) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13243) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6050) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12714) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5610) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20057) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3969) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2272) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21087) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31192) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3987) * $signed(input_fmap_31[7:0]) +
	( 14'sd 8082) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27687) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17805) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22229) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6158) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14840) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18100) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23600) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27298) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8433) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26052) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15458) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26261) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11804) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12054) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23253) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16411) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15725) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24177) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16699) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19139) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29657) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_66[7:0]) +
	( 11'sd 621) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3224) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18595) * $signed(input_fmap_72[7:0]) +
	( 11'sd 715) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4393) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25634) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27945) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12481) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13101) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29623) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14817) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5938) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14372) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7249) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25975) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29127) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7323) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2308) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17252) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32403) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4399) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26919) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15458) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18695) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16067) * $signed(input_fmap_103[7:0]) +
	( 10'sd 275) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9496) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_106[7:0]) +
	( 11'sd 652) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_108[7:0]) +
	( 11'sd 840) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4749) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30489) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29076) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10921) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22578) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19978) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23760) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7448) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17608) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2165) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30353) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5308) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_126[7:0]) +
	( 9'sd 210) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 16'sd 27113) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20054) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21227) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2322) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26060) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27616) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28398) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8590) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7491) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19387) * $signed(input_fmap_16[7:0]) +
	( 11'sd 780) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28076) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29031) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9357) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29862) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7730) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11006) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5597) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5006) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6481) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31164) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15813) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12320) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7254) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9718) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17961) * $signed(input_fmap_40[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23719) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28034) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21348) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28291) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15948) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21766) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1598) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18502) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16338) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15987) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2632) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17658) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9167) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4134) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_61[7:0]) +
	( 10'sd 505) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7494) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29910) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9452) * $signed(input_fmap_68[7:0]) +
	( 9'sd 217) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_70[7:0]) +
	( 11'sd 783) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27642) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3282) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27050) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6946) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3372) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11229) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4594) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10515) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27739) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8517) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23960) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2437) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6526) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27482) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31476) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20268) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7949) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3996) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2572) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9625) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19830) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5185) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22044) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19554) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13053) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4579) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19058) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11866) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23221) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14977) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17081) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2402) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28361) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9547) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21928) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26384) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15518) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30051) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 16'sd 22369) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_3[7:0]) +
	( 13'sd 4038) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11318) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20782) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5786) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28058) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12039) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23926) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9075) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17449) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31052) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18714) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24790) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22876) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18897) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21709) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20056) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14648) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28829) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31121) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31389) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20436) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17166) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10363) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4515) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30105) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2820) * $signed(input_fmap_50[7:0]) +
	( 11'sd 573) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_52[7:0]) +
	( 7'sd 36) * $signed(input_fmap_53[7:0]) +
	( 10'sd 421) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5648) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23396) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10593) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9457) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11465) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17065) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21254) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3115) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24865) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30585) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30025) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29683) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20465) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30062) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28056) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22908) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30895) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21216) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28433) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30761) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16270) * $signed(input_fmap_91[7:0]) +
	( 9'sd 236) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2541) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17436) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_95[7:0]) +
	( 10'sd 272) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22077) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15158) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18693) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12054) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30442) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27649) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11536) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4290) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31570) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16329) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4822) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2314) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4912) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13545) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13934) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2492) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22598) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 15'sd 12877) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18601) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31022) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10913) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26428) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7648) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4217) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18372) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_10[7:0]) +
	( 11'sd 747) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16604) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2473) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16891) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18608) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3754) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13452) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22135) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22944) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29218) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18260) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18207) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1086) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27577) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28677) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17224) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15233) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29502) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13128) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14859) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9777) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1867) * $signed(input_fmap_50[7:0]) +
	( 11'sd 887) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30017) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32314) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18291) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24155) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23510) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8512) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30696) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_64[7:0]) +
	( 13'sd 4044) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31598) * $signed(input_fmap_67[7:0]) +
	( 7'sd 63) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17299) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12659) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31135) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2224) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20959) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_76[7:0]) +
	( 11'sd 526) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7577) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8179) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26710) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5627) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3304) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1086) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9910) * $signed(input_fmap_87[7:0]) +
	( 9'sd 147) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27458) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_90[7:0]) +
	( 10'sd 366) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1676) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16121) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29909) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4683) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5394) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31348) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28016) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26098) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23639) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16023) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16671) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12108) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6051) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26740) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32670) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11260) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13693) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8552) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 16'sd 19671) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6257) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5416) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30099) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7383) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7799) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13376) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9568) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31551) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21492) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31218) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23340) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30726) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28458) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15639) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31661) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26946) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28905) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21857) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25096) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1204) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14921) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22817) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29086) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10639) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27671) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21152) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26297) * $signed(input_fmap_38[7:0]) +
	( 13'sd 4081) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7786) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17142) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21675) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3738) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7400) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21739) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25490) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17896) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22209) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26991) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17477) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7467) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27355) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19896) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19385) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1181) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4543) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29251) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4167) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30432) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7887) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13845) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6785) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29108) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5837) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1033) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10790) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4609) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28793) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26515) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23178) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31582) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17486) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15625) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22921) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21731) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9384) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19226) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14870) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29337) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24517) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19382) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16759) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30734) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25504) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3785) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10951) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30277) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16648) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24771) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30224) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3143) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9143) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10839) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21032) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1718) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30480) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15729) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30738) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5254) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25043) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 16'sd 25903) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17062) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7265) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32296) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25064) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17678) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2704) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22561) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1977) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28519) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24680) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10418) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25321) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26975) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18199) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12790) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20210) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17416) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29237) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14496) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31102) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16510) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25644) * $signed(input_fmap_31[7:0]) +
	( 11'sd 778) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7715) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24730) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29241) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18823) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19746) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_40[7:0]) +
	( 11'sd 634) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5397) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20980) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32316) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28717) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3566) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29220) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2361) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17663) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4286) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6358) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22798) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23552) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6729) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17386) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29611) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2941) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3648) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27929) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6614) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17430) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3480) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14274) * $signed(input_fmap_77[7:0]) +
	( 10'sd 443) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11464) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7171) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6990) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14301) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16532) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14474) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13003) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14631) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20024) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15111) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9531) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28762) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1278) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27378) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30432) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32312) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25589) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27871) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23395) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12204) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29409) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4562) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13384) * $signed(input_fmap_117[7:0]) +
	( 10'sd 370) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10959) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32388) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9098) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 16'sd 17158) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28834) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30080) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14849) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8538) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9173) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11329) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10690) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3544) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3548) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10415) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22031) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30563) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16489) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7812) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15766) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8119) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15085) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20230) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27993) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13531) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6162) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14166) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10534) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29857) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23906) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10825) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4404) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8932) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27549) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15984) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15695) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5545) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14102) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21913) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26502) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12379) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22252) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2497) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9793) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26708) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22551) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20995) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31603) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28719) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31560) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27974) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23623) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28008) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24499) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5533) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21789) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16928) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18618) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29351) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5849) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2572) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19324) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9852) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18902) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12181) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9117) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9358) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4932) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31067) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28425) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27181) * $signed(input_fmap_108[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7652) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24616) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6077) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4409) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9526) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11733) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23050) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5357) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22308) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7467) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 13'sd 2375) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9004) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9367) * $signed(input_fmap_3[7:0]) +
	( 10'sd 375) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18447) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20039) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21484) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16402) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26148) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27490) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21532) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20845) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4721) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20343) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11017) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5254) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25841) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3807) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30790) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1339) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30494) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12131) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9931) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25414) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31893) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_40[7:0]) +
	( 8'sd 113) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23799) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21886) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20514) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23564) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16356) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2160) * $signed(input_fmap_49[7:0]) +
	( 14'sd 8004) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2336) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17663) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6567) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4464) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8742) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7915) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29095) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28341) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17337) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27406) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17681) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24134) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23194) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18921) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_78[7:0]) +
	( 11'sd 736) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13843) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6541) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22742) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8333) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25618) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17333) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10716) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23178) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21626) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20855) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20823) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13888) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8006) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1446) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11575) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2606) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27788) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13427) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30006) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24810) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7498) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23147) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24518) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1800) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28441) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3375) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17189) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_116[7:0]) +
	( 10'sd 506) * $signed(input_fmap_117[7:0]) +
	( 10'sd 358) * $signed(input_fmap_118[7:0]) +
	( 7'sd 45) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22457) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3427) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27112) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5843) * $signed(input_fmap_125[7:0]) +
	( 9'sd 131) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14480) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 16'sd 28325) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5109) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2762) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3881) * $signed(input_fmap_6[7:0]) +
	( 10'sd 495) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11012) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2683) * $signed(input_fmap_9[7:0]) +
	( 10'sd 373) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30678) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14404) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14285) * $signed(input_fmap_14[7:0]) +
	( 11'sd 737) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7309) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31549) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22268) * $signed(input_fmap_19[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_20[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1419) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13364) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8488) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21919) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6106) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26019) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25468) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7696) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8408) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_35[7:0]) +
	( 10'sd 299) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29619) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16029) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5382) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1935) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22002) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16458) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14746) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_52[7:0]) +
	( 11'sd 516) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13732) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20009) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20882) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13646) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11322) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30814) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18161) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23332) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11730) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_71[7:0]) +
	( 11'sd 958) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26909) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5613) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2574) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23293) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2644) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30052) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17196) * $signed(input_fmap_80[7:0]) +
	( 11'sd 970) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25909) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20422) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22982) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31301) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28786) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28411) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6980) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17479) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1681) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13166) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10283) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20877) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32579) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23153) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26593) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32183) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7430) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23818) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8958) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6428) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5388) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31162) * $signed(input_fmap_107[7:0]) +
	( 11'sd 1006) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15362) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22325) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6206) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8260) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18641) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20706) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10550) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16186) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8072) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22309) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 16'sd 22345) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32302) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28937) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1165) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1490) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18660) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27287) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17856) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14631) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15794) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17495) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27887) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26677) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2890) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10703) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7613) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27082) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19043) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17216) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28174) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14317) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17802) * $signed(input_fmap_33[7:0]) +
	( 10'sd 409) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4414) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12333) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23231) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23874) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9588) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13427) * $signed(input_fmap_44[7:0]) +
	( 12'sd 2035) * $signed(input_fmap_45[7:0]) +
	( 4'sd 6) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19905) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29187) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11631) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18545) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2524) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29540) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24912) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1266) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15834) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27729) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26360) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_65[7:0]) +
	( 11'sd 902) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19351) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24830) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8015) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9387) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21497) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1051) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23181) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16489) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26667) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3923) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9188) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24982) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27962) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16935) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30998) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22669) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21852) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32024) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10472) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15631) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21373) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18414) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32205) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19510) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29217) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32540) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6511) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6793) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17662) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27583) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21590) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9689) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29222) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31266) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29719) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20981) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11319) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 13'sd 3031) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13726) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31310) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9102) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18410) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4712) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10358) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22759) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18952) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2484) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32553) * $signed(input_fmap_15[7:0]) +
	( 9'sd 209) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21252) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2555) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19729) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19998) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30882) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32335) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25791) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6901) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22275) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9767) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15386) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9990) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21043) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21191) * $signed(input_fmap_35[7:0]) +
	( 11'sd 684) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3793) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1121) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31428) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2763) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31035) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19103) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17045) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8220) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1952) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32162) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25604) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18239) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3744) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7378) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_60[7:0]) +
	( 11'sd 914) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20170) * $signed(input_fmap_62[7:0]) +
	( 11'sd 957) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5612) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22597) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3389) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20428) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2756) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28137) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4606) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21541) * $signed(input_fmap_74[7:0]) +
	( 10'sd 428) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26565) * $signed(input_fmap_76[7:0]) +
	( 11'sd 542) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17914) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22117) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30674) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4552) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6243) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22663) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29822) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31728) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3467) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25738) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30849) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18261) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29052) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9145) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31687) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16143) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14282) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22838) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2354) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7987) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30089) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6060) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11148) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_117[7:0]) +
	( 11'sd 725) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6768) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32007) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3548) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23108) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4768) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31872) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17534) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13357) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 16'sd 25110) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6237) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_5[7:0]) +
	( 11'sd 886) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27276) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27338) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16697) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24582) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29562) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3001) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23798) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11156) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31856) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15219) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3698) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32209) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29382) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10761) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25558) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22158) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15401) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26635) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18801) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22368) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6337) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11932) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7478) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32466) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32306) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28331) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29533) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26141) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11012) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5251) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8694) * $signed(input_fmap_54[7:0]) +
	( 7'sd 61) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10778) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2666) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12965) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5345) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29779) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30266) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6540) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10014) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3345) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30297) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22731) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4485) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1449) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15160) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1200) * $signed(input_fmap_78[7:0]) +
	( 9'sd 219) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15748) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11856) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31849) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13829) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8800) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11950) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10845) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6230) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30177) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14819) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1332) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14797) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28448) * $signed(input_fmap_100[7:0]) +
	( 10'sd 310) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20620) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3201) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15166) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2652) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5764) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19757) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4648) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29076) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24606) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15848) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22655) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20786) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31482) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27181) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15588) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15775) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21389) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 15'sd 15567) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30077) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10127) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8618) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5230) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2932) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13313) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15624) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18534) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29356) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2906) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5788) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14947) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4900) * $signed(input_fmap_19[7:0]) +
	( 11'sd 781) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9928) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28755) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6307) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2661) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_33[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12987) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6524) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_37[7:0]) +
	( 11'sd 690) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6573) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10737) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23570) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21767) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18653) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25065) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15923) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22828) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3650) * $signed(input_fmap_52[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6384) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28606) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20339) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10173) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32198) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20690) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31094) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5783) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14429) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12858) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9339) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30547) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11183) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15604) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25371) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10535) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12869) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6989) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7342) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8574) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14450) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16062) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24493) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11926) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12266) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18146) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12684) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7706) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2943) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5033) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29280) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5703) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28674) * $signed(input_fmap_102[7:0]) +
	( 11'sd 925) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14197) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22397) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15383) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25882) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25906) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9882) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1754) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14733) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17799) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14396) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9883) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1501) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23203) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25342) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28991) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3735) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24908) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 15'sd 10202) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22834) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12168) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14713) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4225) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24663) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8686) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24739) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26600) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31570) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4325) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32044) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28408) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31018) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_22[7:0]) +
	( 8'sd 97) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11762) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13307) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21321) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1381) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24796) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28494) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28958) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5172) * $signed(input_fmap_36[7:0]) +
	( 11'sd 703) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13418) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3314) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8230) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9321) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24631) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26473) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32358) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6891) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17323) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15723) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12840) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27654) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25707) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16559) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14290) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4222) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5635) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7817) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20424) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30155) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17434) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30294) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31122) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18877) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18081) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2462) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5603) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27337) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20386) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22759) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14622) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3013) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11979) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32355) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9195) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4709) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6924) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15669) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15318) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30056) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8404) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9258) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2322) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14398) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17729) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3347) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26060) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20330) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14364) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5018) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8859) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4465) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15072) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8351) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18824) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26045) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 14'sd 7535) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30787) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5267) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27069) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19793) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17627) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5439) * $signed(input_fmap_10[7:0]) +
	( 11'sd 958) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31782) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24040) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5533) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24022) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6282) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27696) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21822) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11111) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10824) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25441) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12386) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17116) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30625) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7891) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18845) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11896) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3711) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8683) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22305) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11239) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1652) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8243) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20426) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25893) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8208) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9581) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19333) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7740) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19014) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32407) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5942) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28945) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3841) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3789) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9745) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21993) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28716) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20119) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13164) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16926) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11650) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21732) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7915) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28873) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32726) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22055) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5247) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31839) * $signed(input_fmap_82[7:0]) +
	( 11'sd 936) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8920) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3784) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10153) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1261) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30217) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32000) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12240) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7699) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25243) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31538) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11042) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23806) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25835) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14101) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12397) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2915) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2285) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7410) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2381) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19390) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20730) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15575) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16120) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5204) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6662) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3526) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24988) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22636) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 16'sd 31448) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24566) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32502) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26518) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31049) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5381) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26395) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11275) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22998) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13414) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1266) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29362) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24239) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16951) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6435) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3595) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31986) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26187) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18275) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9312) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14919) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26945) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8763) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30022) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26056) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9728) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28037) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11057) * $signed(input_fmap_40[7:0]) +
	( 11'sd 811) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20001) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20946) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22012) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2935) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17318) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20998) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4598) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17946) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29623) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23985) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28671) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30954) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9517) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23414) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27385) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7054) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_64[7:0]) +
	( 11'sd 831) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22352) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10028) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2583) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18032) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11107) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4723) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9575) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30650) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10374) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9162) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3583) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13748) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1254) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18877) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27887) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13278) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32182) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26522) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19395) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1093) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16607) * $signed(input_fmap_95[7:0]) +
	( 11'sd 1001) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11845) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6626) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20877) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9323) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15441) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8072) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23343) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7872) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24084) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31865) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20411) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17494) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15962) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29182) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11519) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18118) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29174) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16375) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32302) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7085) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24865) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7306) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 15'sd 8517) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17623) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18099) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22945) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2628) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1313) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15055) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2246) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1348) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22212) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9415) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19850) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28578) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8664) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5337) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15756) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23522) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28665) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26804) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8615) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27085) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19027) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11730) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23947) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3691) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10135) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19334) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3225) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23174) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22599) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28443) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9793) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8347) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20731) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5266) * $signed(input_fmap_50[7:0]) +
	( 12'sd 2005) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7300) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29371) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16803) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19720) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_57[7:0]) +
	( 11'sd 928) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20092) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18272) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4856) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2149) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32570) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2204) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26369) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25921) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25354) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17516) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1068) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22660) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19181) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14260) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13180) * $signed(input_fmap_86[7:0]) +
	( 9'sd 224) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10877) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21437) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12769) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_95[7:0]) +
	( 11'sd 525) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16692) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29049) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14970) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7133) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7542) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7695) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13607) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9704) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29815) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7211) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17835) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13385) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21784) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13841) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19719) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8657) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13004) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3658) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6247) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28978) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2580) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20387) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19615) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 14'sd 7513) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1159) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30577) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26314) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10388) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21702) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24190) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2429) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11487) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25270) * $signed(input_fmap_14[7:0]) +
	( 14'sd 8031) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16769) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7093) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31440) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31397) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3560) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_25[7:0]) +
	( 11'sd 738) * $signed(input_fmap_26[7:0]) +
	( 9'sd 200) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22025) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23425) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15786) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24954) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3275) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9468) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9326) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5828) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24707) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25159) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1234) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32689) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19478) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11505) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7119) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13177) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3227) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18010) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2855) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11310) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15247) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30548) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22000) * $signed(input_fmap_61[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3686) * $signed(input_fmap_66[7:0]) +
	( 8'sd 125) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21750) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31204) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2148) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17400) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28586) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22610) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15460) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18295) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1761) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_82[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29246) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30540) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23314) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31261) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15449) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24816) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29147) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7979) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22766) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22104) * $signed(input_fmap_98[7:0]) +
	( 11'sd 899) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14598) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18537) * $signed(input_fmap_101[7:0]) +
	( 11'sd 960) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13387) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32156) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19869) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1386) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27979) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17392) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29045) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20556) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26181) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32249) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11632) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27548) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24397) * $signed(input_fmap_121[7:0]) +
	( 10'sd 414) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27974) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5210) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12940) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 13'sd 2561) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18085) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17810) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27958) * $signed(input_fmap_9[7:0]) +
	( 7'sd 35) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3830) * $signed(input_fmap_11[7:0]) +
	( 8'sd 89) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28379) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5247) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10802) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3385) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31490) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19055) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28362) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24493) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2528) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26398) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6440) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27294) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13403) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11240) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10410) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1758) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26241) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1715) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28114) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15470) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18190) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9653) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22744) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31562) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2891) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25485) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12860) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23056) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5843) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18409) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19334) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16865) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3910) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12998) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1995) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4731) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1357) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17452) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31569) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19618) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19064) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10995) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7092) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26986) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18628) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2581) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_92[7:0]) +
	( 7'sd 56) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32555) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13496) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11843) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28328) * $signed(input_fmap_99[7:0]) +
	( 11'sd 647) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22141) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4358) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27820) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30326) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1720) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20712) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3519) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16269) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10740) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27025) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31217) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16679) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16494) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7072) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25868) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 15'sd 14761) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25122) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9353) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16370) * $signed(input_fmap_4[7:0]) +
	( 11'sd 982) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25982) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11636) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9770) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24634) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14487) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18084) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5725) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6299) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31151) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1465) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14973) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2346) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26989) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13711) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21941) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21632) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21515) * $signed(input_fmap_34[7:0]) +
	( 11'sd 875) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10586) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24679) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15506) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6434) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22549) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13266) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29611) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16832) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12446) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25201) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11450) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21116) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10940) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18496) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20107) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19703) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6897) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14175) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11408) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21127) * $signed(input_fmap_70[7:0]) +
	( 12'sd 2012) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2698) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30414) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32281) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8939) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11264) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12027) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30708) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9461) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25458) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9039) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24108) * $signed(input_fmap_93[7:0]) +
	( 10'sd 261) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25498) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31580) * $signed(input_fmap_96[7:0]) +
	( 11'sd 906) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23337) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20004) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9298) * $signed(input_fmap_101[7:0]) +
	( 10'sd 310) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3891) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32554) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11415) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17175) * $signed(input_fmap_112[7:0]) +
	( 10'sd 361) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13822) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_116[7:0]) +
	( 8'sd 108) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_118[7:0]) +
	( 10'sd 390) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23133) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31244) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17448) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30163) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23871) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 16'sd 29693) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25017) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24475) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15137) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6977) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29165) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9600) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1929) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1584) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11549) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5658) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26124) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29521) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8710) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27910) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_26[7:0]) +
	( 11'sd 830) * $signed(input_fmap_27[7:0]) +
	( 11'sd 587) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_30[7:0]) +
	( 9'sd 190) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1425) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12093) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2052) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30349) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1482) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19205) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5062) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25125) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14408) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5849) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28646) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14282) * $signed(input_fmap_48[7:0]) +
	( 11'sd 713) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16382) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8349) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19588) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15819) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10956) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10717) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9389) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6755) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1366) * $signed(input_fmap_60[7:0]) +
	( 8'sd 122) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25727) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12160) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29829) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7954) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10972) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25901) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30038) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3447) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30692) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9700) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12615) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18874) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9250) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12756) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25691) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2116) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22581) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18361) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24390) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3316) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24558) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18448) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3588) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17047) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19377) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13602) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22107) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20224) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8138) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26057) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4828) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28678) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25609) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15597) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22817) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27861) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27875) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25026) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5995) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17467) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25559) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 13'sd 2378) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12689) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13615) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10081) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3071) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12908) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_10[7:0]) +
	( 10'sd 347) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21078) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8366) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29119) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21411) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22967) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8984) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12498) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27818) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2463) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2899) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7792) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9679) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4226) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1552) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15496) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2126) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_42[7:0]) +
	( 11'sd 809) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15877) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2185) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20044) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27278) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30433) * $signed(input_fmap_53[7:0]) +
	( 10'sd 352) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25416) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4803) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31705) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31401) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10257) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22538) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17881) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30823) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22931) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7705) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7478) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29538) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11879) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3839) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18082) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23703) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4378) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16616) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16350) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23679) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18780) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29866) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19021) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7882) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26506) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7368) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27934) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26169) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13264) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10429) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31888) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31469) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6605) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30747) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26565) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8590) * $signed(input_fmap_111[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29483) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_115[7:0]) +
	( 11'sd 855) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15470) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7482) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13446) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32672) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5036) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7966) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20489) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13526) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 16'sd 19753) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9660) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25077) * $signed(input_fmap_2[7:0]) +
	( 11'sd 703) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22786) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31625) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19585) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_8[7:0]) +
	( 8'sd 90) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9347) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20691) * $signed(input_fmap_11[7:0]) +
	( 10'sd 427) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17421) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10736) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3573) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5422) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31630) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24524) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17386) * $signed(input_fmap_23[7:0]) +
	( 11'sd 677) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16441) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17431) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12522) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11843) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9077) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30524) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29189) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32192) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1590) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5367) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24632) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2353) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2829) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24384) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13371) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30244) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25421) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2373) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29736) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20182) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26214) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25957) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9391) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29071) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8870) * $signed(input_fmap_69[7:0]) +
	( 11'sd 513) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6561) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19702) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13566) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10192) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8119) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15002) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31115) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3021) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21728) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11015) * $signed(input_fmap_81[7:0]) +
	( 10'sd 277) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18785) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10421) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16165) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26685) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29214) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26824) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19389) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13809) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8841) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15729) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24980) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24321) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27144) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28522) * $signed(input_fmap_106[7:0]) +
	( 10'sd 381) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25179) * $signed(input_fmap_109[7:0]) +
	( 11'sd 846) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16213) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13759) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_114[7:0]) +
	( 11'sd 535) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23203) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_117[7:0]) +
	( 11'sd 602) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28966) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9028) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15305) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6615) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 16'sd 29334) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9013) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2380) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7042) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23851) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10029) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10180) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24154) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15648) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25764) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18878) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27169) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11633) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5980) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8222) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30222) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27033) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24506) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12466) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5484) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17535) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18627) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23262) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14547) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18492) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8524) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13311) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26699) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13073) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27500) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29469) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25444) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17602) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7341) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28164) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20352) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22456) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14056) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6385) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7295) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1892) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20618) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1106) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5528) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_58[7:0]) +
	( 6'sd 27) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15764) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2494) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29037) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14901) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1829) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21754) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9026) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22974) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21326) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21397) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24584) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22229) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11095) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11734) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3378) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8595) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9009) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19277) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23680) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14905) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21655) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10535) * $signed(input_fmap_91[7:0]) +
	( 10'sd 309) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6569) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25375) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8556) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21912) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26103) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3474) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8854) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19224) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31298) * $signed(input_fmap_117[7:0]) +
	( 7'sd 47) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17268) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24887) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23503) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27615) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11093) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 16'sd 19208) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13462) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19623) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29423) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4391) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26047) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8558) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10510) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26199) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2874) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23208) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2920) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29678) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15931) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22964) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26387) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11185) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31597) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20068) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6759) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21309) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8113) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12268) * $signed(input_fmap_38[7:0]) +
	( 10'sd 494) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2692) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23764) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3622) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26271) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32479) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21193) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23231) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18551) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32307) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8253) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21597) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25844) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22036) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25574) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_66[7:0]) +
	( 11'sd 577) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12191) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21109) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23100) * $signed(input_fmap_74[7:0]) +
	( 11'sd 572) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9518) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4919) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13739) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18726) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28157) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11066) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22737) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30114) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27789) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1667) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32572) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24113) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15480) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5808) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28698) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8481) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19968) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9867) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16396) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_110[7:0]) +
	( 11'sd 611) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27989) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18050) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8574) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21579) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23001) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10271) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18776) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32729) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6889) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14878) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 15'sd 9233) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27126) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20298) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5218) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30337) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16010) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23559) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3415) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27454) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13211) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10520) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3055) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18081) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24079) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30115) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18279) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16339) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12828) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15441) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14164) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27326) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15925) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27101) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13700) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32545) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5405) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20787) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32598) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13144) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11334) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18041) * $signed(input_fmap_46[7:0]) +
	( 11'sd 730) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28655) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3405) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14970) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13371) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19538) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9865) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10273) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24274) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29311) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22510) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14361) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20687) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10076) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1230) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27868) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31622) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14873) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22262) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16792) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29893) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22228) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26917) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6245) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15643) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3846) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_91[7:0]) +
	( 10'sd 504) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25924) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18605) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20828) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23288) * $signed(input_fmap_98[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3378) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8972) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15921) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24632) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17084) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5921) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9779) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1152) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25097) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30811) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23551) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24603) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21491) * $signed(input_fmap_118[7:0]) +
	( 11'sd 667) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27155) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9085) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19003) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19050) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10585) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21842) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 15'sd 9762) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15903) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14919) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27458) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_5[7:0]) +
	( 11'sd 763) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12108) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8970) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6605) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19560) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1800) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7964) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32161) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6132) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8829) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26295) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3560) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6420) * $signed(input_fmap_30[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_31[7:0]) +
	( 13'sd 4053) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4383) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9684) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3840) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31798) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13159) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25655) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14313) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2978) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30665) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25689) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26725) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30529) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16440) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10005) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5123) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2292) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4592) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16017) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3622) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16760) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19643) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26774) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1825) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3024) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8641) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16792) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28209) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23041) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22942) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21009) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15946) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27950) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21375) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7050) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31442) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13849) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14171) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23106) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7388) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7412) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8041) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27870) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23579) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29535) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16968) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17953) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32448) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17483) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22380) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14606) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20457) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3379) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6166) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23387) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19640) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13444) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18199) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27925) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20583) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 15'sd 12595) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10929) * $signed(input_fmap_1[7:0]) +
	( 13'sd 4090) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32495) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3504) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12178) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20182) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21676) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7238) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27603) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20331) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25329) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31612) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21097) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13385) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31150) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_17[7:0]) +
	( 12'sd 2018) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10703) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7399) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10279) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6897) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21209) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29852) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17373) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10342) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24562) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15772) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11976) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19904) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17852) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23848) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27564) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12714) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16545) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_46[7:0]) +
	( 11'sd 908) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11357) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8521) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23250) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16749) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11977) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16989) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10921) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27554) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32521) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2107) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31776) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10656) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11386) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8655) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4530) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14436) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25673) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1895) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28774) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22633) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18166) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26343) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3281) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24473) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7439) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_80[7:0]) +
	( 11'sd 664) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14153) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9449) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27273) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21663) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7098) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29720) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30040) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12431) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11795) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30134) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27224) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19440) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27772) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23297) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16050) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17937) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11391) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14015) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20987) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19667) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11768) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30938) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26493) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19997) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12835) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28593) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9095) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19643) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12594) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16844) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_119[7:0]) +
	( 11'sd 656) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2821) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_123[7:0]) +
	( 11'sd 684) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17815) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24948) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22336) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 14'sd 5364) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29576) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7225) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_4[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7664) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32341) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25744) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31824) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28568) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28626) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23872) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17988) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24397) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14313) * $signed(input_fmap_21[7:0]) +
	( 11'sd 720) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27564) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30707) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20323) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5324) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4326) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27510) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25908) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19971) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12518) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3823) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4582) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21399) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6423) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4168) * $signed(input_fmap_42[7:0]) +
	( 11'sd 680) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32636) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29699) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17279) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10005) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32093) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25704) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16924) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5798) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7428) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6325) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8091) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14983) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15715) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20712) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1849) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19694) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5242) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20514) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1948) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14851) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28751) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24683) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18594) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_78[7:0]) +
	( 13'sd 4016) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24729) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29533) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29880) * $signed(input_fmap_84[7:0]) +
	( 11'sd 529) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5744) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20328) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18602) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4920) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3424) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6924) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23170) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31234) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31654) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19288) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18560) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7952) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16408) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30292) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11234) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18897) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30069) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12999) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12114) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14966) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25782) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21389) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28102) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 16'sd 28805) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6325) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8964) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18765) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18469) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15830) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25883) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15614) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11003) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13214) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28981) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18910) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3989) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13882) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32418) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28795) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27621) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5879) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17458) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20660) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_32[7:0]) +
	( 12'sd 2030) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13490) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10742) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22304) * $signed(input_fmap_36[7:0]) +
	( 11'sd 611) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9142) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30152) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15201) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_42[7:0]) +
	( 11'sd 740) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14851) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19729) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1674) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17546) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7577) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9794) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15101) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13845) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18973) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2917) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23819) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22705) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22328) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15173) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7034) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12596) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8294) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23295) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15964) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23646) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20176) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13189) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7473) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13371) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16893) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12759) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6979) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5382) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18403) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2122) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6768) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26361) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5962) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15181) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30411) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3197) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26206) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7841) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19265) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29416) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12214) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21064) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11037) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21712) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31735) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22185) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15873) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11358) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2219) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23837) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14024) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23761) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14947) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28764) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30698) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27611) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 16'sd 17095) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30745) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14856) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26689) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16162) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31860) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21713) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20141) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16104) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21070) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29094) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32713) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12134) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2677) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2597) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24488) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19724) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28469) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16807) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18945) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4566) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2957) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18669) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15397) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18576) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14770) * $signed(input_fmap_42[7:0]) +
	( 11'sd 881) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11181) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24410) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31288) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1339) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3816) * $signed(input_fmap_50[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6952) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11011) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23250) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21963) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10604) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17579) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3409) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29903) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6631) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6413) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8249) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6358) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26781) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23989) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10071) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14057) * $signed(input_fmap_73[7:0]) +
	( 11'sd 757) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12483) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26601) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14908) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25636) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19172) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32394) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21920) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31442) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28359) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12967) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7165) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31239) * $signed(input_fmap_97[7:0]) +
	( 8'sd 126) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13247) * $signed(input_fmap_100[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6498) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21804) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15971) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10415) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5510) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30890) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25769) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16979) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17891) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22354) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32425) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12163) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 14'sd 7583) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7419) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10516) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5040) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30151) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10214) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6141) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31552) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14935) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27963) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19445) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10968) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6664) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29909) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6396) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16802) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7602) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20282) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11343) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30603) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20810) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24249) * $signed(input_fmap_33[7:0]) +
	( 14'sd 8040) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23846) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21848) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21285) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22077) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30725) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24575) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31975) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24157) * $signed(input_fmap_44[7:0]) +
	( 11'sd 981) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26914) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24751) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21276) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4439) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23766) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9323) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25999) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3280) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16840) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25391) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7287) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15099) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15966) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22031) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25270) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19783) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6480) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9583) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27354) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5618) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28025) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_77[7:0]) +
	( 9'sd 140) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31586) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5592) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27212) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7680) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24701) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19491) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9189) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23976) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10542) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8281) * $signed(input_fmap_98[7:0]) +
	( 11'sd 525) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17717) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10333) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1479) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14950) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3451) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6664) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3308) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32713) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15397) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18656) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10392) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11630) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28999) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18983) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29241) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12877) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8888) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 16'sd 17849) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22317) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13485) * $signed(input_fmap_2[7:0]) +
	( 8'sd 94) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7629) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4289) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2559) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16180) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_9[7:0]) +
	( 11'sd 635) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16659) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9115) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21962) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7019) * $signed(input_fmap_16[7:0]) +
	( 14'sd 8124) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12355) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9107) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20979) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21661) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20823) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8865) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5123) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31275) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26083) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29140) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9174) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9108) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10258) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3537) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9111) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32563) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15446) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11241) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10461) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13364) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30870) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8512) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30860) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20785) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12521) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26202) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22711) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4547) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31028) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18178) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7759) * $signed(input_fmap_72[7:0]) +
	( 13'sd 4071) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9437) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13056) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26278) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13248) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18061) * $signed(input_fmap_79[7:0]) +
	( 13'sd 4071) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16076) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9732) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24106) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31955) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7075) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27545) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18166) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24973) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7160) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16516) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20706) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10717) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19180) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12702) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2296) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23848) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23725) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4256) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21416) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5902) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22463) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3099) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19405) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20378) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32194) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3607) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15715) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32645) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16277) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2355) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19556) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12906) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24124) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15453) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 12'sd 1286) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26490) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_3[7:0]) +
	( 14'sd 8127) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13780) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11303) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19305) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23102) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19970) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17353) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16588) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9603) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22887) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15323) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8221) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21292) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30344) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6306) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21021) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10408) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10461) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3417) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6318) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30940) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8961) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3671) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14009) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26257) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5255) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17370) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5158) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15096) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4716) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12820) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6843) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8481) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1128) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4600) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4638) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6127) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15474) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2919) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27108) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18123) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14346) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4128) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25864) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6813) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3835) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13708) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26515) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25287) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7240) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27820) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32064) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16371) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13820) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3970) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21235) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3085) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14293) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28740) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25519) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12042) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9333) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32546) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21352) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25908) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2442) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_124[7:0]) +
	( 5'sd 12) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14818) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 16'sd 19250) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4617) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12324) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23833) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14631) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16648) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24503) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11377) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17406) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10698) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18696) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3915) * $signed(input_fmap_17[7:0]) +
	( 11'sd 701) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3870) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13981) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24678) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9337) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27347) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12326) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30370) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4188) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17101) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21043) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21093) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3047) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11571) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15106) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16724) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26593) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4487) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25567) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32761) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28950) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_53[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1071) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11585) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10980) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8996) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21699) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15492) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12636) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10832) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23769) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25973) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7162) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17863) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24932) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31586) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25696) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29440) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14061) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29845) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9952) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28146) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15583) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14791) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19800) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20665) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7106) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2531) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31046) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12084) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3715) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17440) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11880) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7922) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16314) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25125) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2619) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18396) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31968) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18295) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20115) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12214) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3632) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22955) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29829) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5410) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8268) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13071) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_114[7:0]) +
	( 10'sd 388) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23426) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30280) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26746) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6921) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3731) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20744) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12324) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19151) * $signed(input_fmap_125[7:0]) +
	( 10'sd 258) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5250) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 16'sd 28624) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19851) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32617) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30435) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17944) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17555) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22802) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7259) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17658) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12892) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7278) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2055) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24144) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22243) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9045) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29249) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28759) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1692) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31307) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31780) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3309) * $signed(input_fmap_32[7:0]) +
	( 10'sd 390) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7994) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12891) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24606) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4114) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3876) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7529) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32314) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15722) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23088) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17506) * $signed(input_fmap_53[7:0]) +
	( 11'sd 795) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8528) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22942) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4118) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15914) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23643) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14480) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28937) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4397) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12696) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7895) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14061) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27576) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29379) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21742) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1077) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12932) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18994) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4949) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4579) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5011) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24612) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17602) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29733) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12358) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22278) * $signed(input_fmap_91[7:0]) +
	( 11'sd 623) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6908) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9349) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7871) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18933) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8660) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16371) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23300) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9485) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5804) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21101) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10810) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9842) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24797) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25485) * $signed(input_fmap_121[7:0]) +
	( 9'sd 200) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32528) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17147) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19101) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 16'sd 24688) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23175) * $signed(input_fmap_1[7:0]) +
	( 11'sd 523) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19407) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22277) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18716) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4807) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31376) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6866) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11171) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26539) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19196) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4373) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22232) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27020) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23821) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25849) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6316) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10942) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16797) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20706) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29072) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31369) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8250) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2680) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17318) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11708) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11473) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17919) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16733) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22973) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11246) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2235) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11128) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10806) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15754) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14053) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5494) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27347) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31666) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16591) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27044) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26739) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20973) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26891) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6340) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28773) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11830) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22690) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12965) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18444) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12125) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24497) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24817) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30773) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5394) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18174) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25759) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20909) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21619) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30297) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12585) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6245) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30180) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7853) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8752) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8543) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30488) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8694) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17487) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27738) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19771) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4219) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27761) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27213) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1631) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32176) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26296) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2923) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12596) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4371) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14201) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9366) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12902) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30911) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30690) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21141) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25056) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 14'sd 5153) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20701) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23771) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6098) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3208) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28141) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25439) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3960) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2085) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5809) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16181) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4219) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1736) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12919) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4921) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19065) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7466) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26817) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10441) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21877) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9647) * $signed(input_fmap_30[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12909) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25173) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31402) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14874) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12976) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32014) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25421) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11143) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15944) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3255) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29836) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5320) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24735) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18676) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14045) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21655) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13593) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_57[7:0]) +
	( 7'sd 43) * $signed(input_fmap_58[7:0]) +
	( 8'sd 105) * $signed(input_fmap_59[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23476) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25492) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6948) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29646) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19145) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1997) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3319) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11179) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20810) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6307) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20948) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_83[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9912) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28314) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8233) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14904) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19720) * $signed(input_fmap_93[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4396) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20797) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22256) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1215) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27958) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10927) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32030) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4342) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14053) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28347) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16184) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19040) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7436) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13289) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13616) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8678) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31526) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18311) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24536) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6651) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5388) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21420) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28336) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 16'sd 28908) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_2[7:0]) +
	( 12'sd 2014) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28448) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6648) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19600) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20798) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13226) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12845) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2092) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31116) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20137) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11610) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32329) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20352) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18883) * $signed(input_fmap_24[7:0]) +
	( 11'sd 905) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31653) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11422) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12565) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23176) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14768) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26334) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21008) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24957) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3555) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26862) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30098) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22115) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12158) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27303) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32535) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15762) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27446) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23815) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24854) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21879) * $signed(input_fmap_49[7:0]) +
	( 11'sd 524) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2219) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13343) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8309) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6409) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_59[7:0]) +
	( 9'sd 148) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31396) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23931) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24486) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6292) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14440) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12639) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27220) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9417) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19247) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1366) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16212) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26812) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6587) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18250) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12882) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10609) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4693) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14150) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7831) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12158) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30813) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24225) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28055) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11618) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2672) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4856) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4345) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22397) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18676) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5403) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24770) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28331) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8596) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10197) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31365) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28938) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23442) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5047) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7328) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25128) * $signed(input_fmap_126[7:0]) +
	( 8'sd 103) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 18229) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5406) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24989) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17553) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19355) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18483) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16302) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9802) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26369) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29260) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4188) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10398) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27868) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3287) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1905) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27057) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28643) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12818) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1575) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3734) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23526) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16461) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29945) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21914) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4391) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32380) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17125) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15516) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11299) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20789) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9379) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32162) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3961) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16599) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28501) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2700) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24650) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26412) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16489) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16876) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32215) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25755) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11798) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16225) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23483) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31053) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9088) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1789) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4140) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25506) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26056) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23195) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18504) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27798) * $signed(input_fmap_93[7:0]) +
	( 14'sd 8185) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14063) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3029) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_98[7:0]) +
	( 11'sd 983) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18605) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25974) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3032) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28882) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9423) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26955) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3754) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15360) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12754) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10335) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12899) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3677) * $signed(input_fmap_119[7:0]) +
	( 11'sd 607) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4889) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21807) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9236) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2637) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 14'sd 7119) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21975) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5221) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15300) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6344) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22262) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21424) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27287) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10732) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16629) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12293) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9322) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2973) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14361) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9730) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15984) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26711) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28261) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5749) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20478) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3098) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9653) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6995) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9608) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14123) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16734) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17416) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24922) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10293) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1695) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26714) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29923) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29488) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25204) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1823) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22807) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19871) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13687) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3904) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29278) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25290) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10032) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14355) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13345) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5346) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23731) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10347) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28963) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6992) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13798) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24453) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26934) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14571) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10938) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19691) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7903) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24807) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18492) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30163) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30685) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12954) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24713) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11331) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25894) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4250) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26576) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15178) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9942) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27939) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18617) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7732) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2767) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15363) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31050) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31701) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21137) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18914) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30907) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16408) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1527) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 16'sd 19064) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7617) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2538) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21225) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8963) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8715) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6772) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25279) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19347) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13454) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27884) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9988) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2968) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30259) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12063) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25062) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30899) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20739) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2822) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11021) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2981) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14463) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31420) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21204) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31688) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29234) * $signed(input_fmap_48[7:0]) +
	( 11'sd 651) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30650) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7694) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12758) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15233) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_58[7:0]) +
	( 11'sd 884) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11704) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1620) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6849) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12764) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14699) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30279) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1325) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3967) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8663) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27753) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6674) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6804) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4817) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1606) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4184) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29021) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24770) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_85[7:0]) +
	( 11'sd 596) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9492) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26840) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19726) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_93[7:0]) +
	( 11'sd 611) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12312) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6516) * $signed(input_fmap_99[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19451) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8871) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27184) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28045) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21225) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12096) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17537) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3963) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28254) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21418) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31749) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17578) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30748) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7549) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31812) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_119[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11589) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32757) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13843) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12924) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13512) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 15'sd 13446) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16135) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15372) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31775) * $signed(input_fmap_5[7:0]) +
	( 10'sd 432) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22840) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14669) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30746) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5142) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_15[7:0]) +
	( 11'sd 585) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4397) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28008) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15793) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22645) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25424) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28528) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8970) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29690) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8626) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_29[7:0]) +
	( 11'sd 570) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20665) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19497) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31736) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24947) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21549) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10319) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7445) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12796) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29694) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22434) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18193) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4241) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7058) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16810) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23299) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2699) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19691) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30792) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10351) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7179) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3375) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20815) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2954) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25966) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12569) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24197) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21458) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14599) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6694) * $signed(input_fmap_75[7:0]) +
	( 10'sd 295) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11719) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22506) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25964) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21486) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20574) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8457) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3956) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2544) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9454) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1657) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10782) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5864) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23778) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14556) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27332) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29987) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32018) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20344) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30906) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12225) * $signed(input_fmap_104[7:0]) +
	( 8'sd 103) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24137) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28292) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10791) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13849) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15454) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26634) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5881) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30521) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26156) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15249) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21874) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18143) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15341) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24250) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 15'sd 12064) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17906) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14396) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20611) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9251) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22393) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26039) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25359) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15129) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20575) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11189) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23917) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30864) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6911) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29075) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18837) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10453) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32730) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2539) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23402) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31106) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5672) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25419) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28711) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19463) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30650) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3345) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25605) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24298) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26461) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30442) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2938) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24017) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14365) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21353) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13348) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25999) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5675) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26116) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23013) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27883) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21009) * $signed(input_fmap_71[7:0]) +
	( 7'sd 62) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28306) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20973) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4769) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28756) * $signed(input_fmap_77[7:0]) +
	( 10'sd 495) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29396) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1853) * $signed(input_fmap_80[7:0]) +
	( 9'sd 146) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24711) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20269) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31545) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24052) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18843) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5388) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12809) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12875) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2638) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27305) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1282) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30253) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5221) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24387) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10442) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17146) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7013) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9802) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11170) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25920) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15997) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17551) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7662) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3592) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17947) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12691) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17389) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22167) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 13'sd 3681) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27941) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3782) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19045) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5067) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18115) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32493) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3341) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16602) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5426) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17043) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7322) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12843) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21568) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13953) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30882) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16361) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10696) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25573) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12751) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25751) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17542) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16073) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15291) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10366) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26892) * $signed(input_fmap_37[7:0]) +
	( 8'sd 122) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15621) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24685) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16114) * $signed(input_fmap_43[7:0]) +
	( 8'sd 115) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18996) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10403) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16513) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23185) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2328) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22110) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30634) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22601) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29578) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6438) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29719) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1708) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13852) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28187) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16269) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9891) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6341) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21654) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5248) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25301) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6093) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32489) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20457) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13906) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23523) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25774) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12921) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20188) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31149) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26795) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25296) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5384) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17113) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14106) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18622) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24165) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17572) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20441) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13033) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19899) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13073) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19186) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13243) * $signed(input_fmap_112[7:0]) +
	( 11'sd 879) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13564) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19085) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23133) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24678) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6262) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22839) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14585) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8854) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30656) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17847) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24700) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 13'sd 3597) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20171) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13149) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27070) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18856) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23337) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28226) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3051) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20439) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13746) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7795) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2462) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28198) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2771) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27415) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20713) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22300) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23116) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4932) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15078) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10286) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23263) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29985) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10118) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16735) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21365) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5293) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13211) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16362) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9298) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25845) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31226) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_54[7:0]) +
	( 11'sd 578) * $signed(input_fmap_55[7:0]) +
	( 11'sd 882) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19972) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24832) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17471) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11146) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8306) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13919) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12050) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18590) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16214) * $signed(input_fmap_67[7:0]) +
	( 10'sd 415) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22507) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1337) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2632) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18656) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25254) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7120) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9534) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10498) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1069) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22446) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7942) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2951) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2669) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7517) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1129) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27477) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25452) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18796) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18186) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3265) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18570) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12232) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9550) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13265) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29894) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2224) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19106) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10395) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18457) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10249) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3674) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16919) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16414) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14705) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25718) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21842) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28463) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3401) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30930) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21840) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14051) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24534) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 15'sd 13378) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29142) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28120) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13729) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28579) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3327) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26086) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20202) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8762) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21562) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11130) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24950) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8733) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32132) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1415) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20791) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3854) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5321) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9828) * $signed(input_fmap_33[7:0]) +
	( 9'sd 216) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24792) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18373) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6025) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23967) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21004) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2871) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19066) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32141) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12791) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27993) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16336) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8211) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8759) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_53[7:0]) +
	( 8'sd 95) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24839) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24594) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16775) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12009) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31213) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4920) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24635) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4849) * $signed(input_fmap_63[7:0]) +
	( 11'sd 909) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4195) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27506) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23278) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31698) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31558) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26976) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_78[7:0]) +
	( 9'sd 149) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24604) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4617) * $signed(input_fmap_82[7:0]) +
	( 6'sd 23) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9043) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8531) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30940) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19049) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19573) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20640) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5891) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25458) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30758) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16007) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24905) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6412) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4492) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20934) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12116) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17841) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4571) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3385) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26662) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17252) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25028) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20294) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9376) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9515) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27402) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23386) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23137) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9807) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9380) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27791) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8231) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 12'sd 1855) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30486) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11356) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10916) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5163) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6467) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3567) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4636) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10665) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7108) * $signed(input_fmap_11[7:0]) +
	( 10'sd 462) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11331) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8574) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10894) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19506) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1441) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17387) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31349) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3604) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10425) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16076) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11124) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21616) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5366) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26653) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28764) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4900) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18119) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31273) * $signed(input_fmap_42[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18561) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31190) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6378) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4483) * $signed(input_fmap_62[7:0]) +
	( 10'sd 470) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8588) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13324) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19626) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12801) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30276) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29267) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24855) * $signed(input_fmap_74[7:0]) +
	( 14'sd 8090) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18660) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20889) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23172) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11578) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14797) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21857) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30418) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6631) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32371) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32021) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4102) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21051) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30072) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9911) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6341) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29210) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25515) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21402) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25438) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12738) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15001) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12137) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3293) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16752) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3426) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5079) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21975) * $signed(input_fmap_120[7:0]) +
	( 8'sd 83) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22238) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10548) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22004) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 16'sd 25046) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20960) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6811) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9415) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4217) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15017) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23579) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16724) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26640) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4910) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26353) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6159) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24479) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22993) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20658) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18448) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23710) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6591) * $signed(input_fmap_30[7:0]) +
	( 9'sd 223) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6542) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_36[7:0]) +
	( 10'sd 468) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7941) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23082) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21724) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15344) * $signed(input_fmap_43[7:0]) +
	( 11'sd 804) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8768) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12235) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3816) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21874) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12691) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9449) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29353) * $signed(input_fmap_59[7:0]) +
	( 9'sd 148) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1343) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7298) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13069) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4473) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19455) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18425) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1753) * $signed(input_fmap_72[7:0]) +
	( 13'sd 4086) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20836) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21934) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29850) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4369) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5650) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16128) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18863) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23957) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8911) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12842) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4286) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19083) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29562) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20170) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30830) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2629) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23644) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10010) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16326) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2533) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4828) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19866) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7646) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18650) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25850) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19418) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13086) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13005) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3524) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15225) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25005) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14361) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17361) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13433) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30012) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30620) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 16'sd 26146) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17015) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21437) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30382) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16798) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7279) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28041) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23815) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5242) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17253) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18935) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11215) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13591) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28539) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30978) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3845) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27183) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5837) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25689) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2357) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16622) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17993) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13878) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28081) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24618) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29796) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28739) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25401) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4900) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8570) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4431) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2788) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8134) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24300) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19758) * $signed(input_fmap_55[7:0]) +
	( 10'sd 390) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4997) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7290) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26921) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31085) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4534) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30956) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17261) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2639) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9866) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25252) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18490) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11727) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16725) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3231) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9120) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26516) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31062) * $signed(input_fmap_78[7:0]) +
	( 11'sd 937) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6385) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_84[7:0]) +
	( 11'sd 799) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30203) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1900) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13680) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28524) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6869) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7306) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29761) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23652) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3287) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15143) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6219) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20925) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23863) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31072) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2349) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24525) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21513) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26052) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3190) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30355) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21924) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 16'sd 21817) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8818) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26867) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28766) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5734) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15519) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23921) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17134) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8140) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21493) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12548) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16457) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22397) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6337) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6706) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23960) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14933) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17908) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2383) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1556) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2943) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_30[7:0]) +
	( 13'sd 4056) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29474) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31795) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4624) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2207) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25212) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31718) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11749) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21586) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23638) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21928) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23698) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1860) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24155) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15418) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5170) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14401) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15324) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23011) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10825) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25726) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13468) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3990) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30590) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17612) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3087) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24849) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32302) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8908) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9783) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23109) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20725) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6353) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32467) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7310) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13362) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14163) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28239) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23324) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1255) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27293) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9813) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21883) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9112) * $signed(input_fmap_105[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13827) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31071) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17161) * $signed(input_fmap_110[7:0]) +
	( 7'sd 40) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16669) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18474) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6229) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4411) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30422) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19047) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1691) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9539) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_123[7:0]) +
	( 11'sd 585) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28591) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6907) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 12'sd 1815) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26741) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28179) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16254) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15937) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2985) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11788) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18400) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2843) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16964) * $signed(input_fmap_17[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27183) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25134) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7541) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15733) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30386) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5058) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15568) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26775) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21459) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25678) * $signed(input_fmap_31[7:0]) +
	( 11'sd 734) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15578) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8721) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19844) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31821) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21233) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5191) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12288) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29644) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4481) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15159) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13384) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15107) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7696) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24965) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26059) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29420) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25171) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29943) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11867) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1524) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17402) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11838) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18604) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_74[7:0]) +
	( 10'sd 292) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26250) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1440) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30328) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1606) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6845) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14775) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17581) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23606) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20865) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28588) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10005) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26516) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22460) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17794) * $signed(input_fmap_102[7:0]) +
	( 11'sd 707) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28709) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17139) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24702) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18332) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_113[7:0]) +
	( 11'sd 553) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2333) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16211) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29511) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4497) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16538) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28634) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3886) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4263) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2150) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10470) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6679) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 16'sd 26903) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13691) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21263) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7902) * $signed(input_fmap_3[7:0]) +
	( 7'sd 57) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28905) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23210) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29448) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32528) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13777) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32008) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21694) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28593) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3635) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21268) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9344) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16123) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20298) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28727) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27904) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20165) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32340) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4511) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4941) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30743) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29275) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30544) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24383) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22874) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16092) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10982) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22779) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26000) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12450) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12893) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4466) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29591) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_51[7:0]) +
	( 10'sd 397) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1437) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31821) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5064) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20617) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4658) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27413) * $signed(input_fmap_65[7:0]) +
	( 9'sd 196) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3387) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6078) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2971) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_71[7:0]) +
	( 10'sd 270) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21280) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8837) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8139) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1963) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29521) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5468) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1206) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22404) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28157) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21831) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25968) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10289) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31790) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16205) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26959) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4114) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19140) * $signed(input_fmap_97[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15873) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29412) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19591) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13289) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28770) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21298) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5152) * $signed(input_fmap_111[7:0]) +
	( 14'sd 8080) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31016) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21874) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12820) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6650) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16981) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31541) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23384) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22043) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15693) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5164) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6054) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 14'sd 4735) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15050) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11269) * $signed(input_fmap_3[7:0]) +
	( 11'sd 746) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1464) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3155) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11652) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21864) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18302) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15690) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18506) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21260) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5052) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2990) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28720) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6781) * $signed(input_fmap_22[7:0]) +
	( 11'sd 512) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18162) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2874) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32472) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20618) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6619) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25252) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3383) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11074) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31246) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28906) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10329) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7203) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7840) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26254) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2909) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_47[7:0]) +
	( 11'sd 659) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6677) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15267) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18284) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10113) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24105) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17832) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21303) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29290) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3092) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6012) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8517) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23934) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3316) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26194) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16497) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11306) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9216) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4689) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22912) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17641) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29494) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20715) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15202) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20503) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28952) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12969) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9168) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29230) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22672) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31694) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5459) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5865) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4447) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7459) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25649) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12617) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6617) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20295) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17563) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_109[7:0]) +
	( 10'sd 350) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26351) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31037) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15553) * $signed(input_fmap_115[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14175) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26570) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1366) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14354) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24706) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7151) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10677) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 16'sd 19296) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10071) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19649) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29470) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29326) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18723) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4382) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22682) * $signed(input_fmap_9[7:0]) +
	( 11'sd 592) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20997) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9632) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23202) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26197) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3087) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15883) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18774) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31445) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27958) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31177) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12710) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20920) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20167) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24163) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13120) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15878) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12800) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10379) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5140) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25442) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_46[7:0]) +
	( 12'sd 2034) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3397) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23752) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27486) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17448) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23155) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21175) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13894) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18638) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17735) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24793) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16468) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25677) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25465) * $signed(input_fmap_65[7:0]) +
	( 7'sd 51) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8973) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31545) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25574) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25555) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9932) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15407) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_75[7:0]) +
	( 11'sd 711) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4657) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2161) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22258) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24371) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14017) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11726) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2255) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13185) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32343) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1690) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13819) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17244) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18996) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29762) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2330) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27815) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9731) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8499) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26553) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29226) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11899) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17808) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12595) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3748) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22102) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25599) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3329) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_125[7:0]) +
	( 14'sd 8029) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19243) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 14'sd 5038) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10837) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13287) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1130) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7266) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19086) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4402) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30202) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24453) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_26[7:0]) +
	( 11'sd 701) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25315) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28247) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9517) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14149) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27389) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19617) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21524) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18111) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15034) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27556) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7025) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25176) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16356) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30566) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11061) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14178) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18340) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21620) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12803) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29232) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14333) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32410) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6030) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20437) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4271) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17166) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28266) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9608) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7814) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12426) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15098) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25536) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16734) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25297) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25930) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25251) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16474) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23789) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2988) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6584) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23274) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27170) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29510) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5049) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6114) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11578) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12161) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26836) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16909) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27677) * $signed(input_fmap_102[7:0]) +
	( 8'sd 81) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10825) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32336) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_106[7:0]) +
	( 8'sd 82) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15385) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2941) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23593) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14101) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12396) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18437) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2191) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21853) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20151) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20265) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31582) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15476) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_125[7:0]) +
	( 10'sd 349) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 15'sd 11065) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20513) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10996) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12492) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12042) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_11[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16532) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5689) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_15[7:0]) +
	( 10'sd 473) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29840) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23622) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14296) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20050) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3807) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4770) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13325) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20448) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2284) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29488) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24511) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20617) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11488) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2638) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10922) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25887) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7841) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21501) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31216) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1833) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18064) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30078) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15917) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25488) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8768) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18250) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29293) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10659) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20094) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13924) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17636) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26754) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6769) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19434) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16160) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11292) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8344) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24461) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20084) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23464) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21420) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32167) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30557) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18089) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7935) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19727) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20246) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15012) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25769) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23035) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29272) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19372) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4376) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14308) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4760) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18337) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6191) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20504) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2495) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14295) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17857) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23001) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18595) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29452) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9043) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22115) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26347) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28638) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18094) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17910) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11759) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 15'sd 8711) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20045) * $signed(input_fmap_4[7:0]) +
	( 11'sd 517) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21712) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7579) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1721) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5139) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7267) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31595) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8199) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13033) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12351) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5181) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14717) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26508) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14687) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4556) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29579) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9353) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30281) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29524) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11390) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32090) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29464) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3418) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24085) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2691) * $signed(input_fmap_50[7:0]) +
	( 6'sd 21) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5423) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11471) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27653) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17550) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10236) * $signed(input_fmap_67[7:0]) +
	( 14'sd 8076) * $signed(input_fmap_68[7:0]) +
	( 11'sd 676) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18536) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20150) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1705) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25940) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21102) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8548) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5881) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5597) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9256) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31169) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25495) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19779) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7338) * $signed(input_fmap_86[7:0]) +
	( 5'sd 10) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4893) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7972) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6565) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16673) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22866) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24512) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16138) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17223) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21937) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21267) * $signed(input_fmap_100[7:0]) +
	( 11'sd 868) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20374) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24524) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18989) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17406) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19844) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3113) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13275) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13844) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30384) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7721) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10471) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7466) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2951) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24976) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7278) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4355) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14796) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 12'sd 1469) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3532) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25677) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24642) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16657) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27166) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9078) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9204) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14309) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9667) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22885) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4111) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3269) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13346) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2349) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22510) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30981) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31905) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15822) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27926) * $signed(input_fmap_37[7:0]) +
	( 10'sd 367) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18782) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26561) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21252) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32483) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9738) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2055) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1253) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7446) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16293) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9117) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25503) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14403) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30936) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18253) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25153) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27967) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13917) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9007) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16145) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24488) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4848) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32059) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13774) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21006) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21264) * $signed(input_fmap_73[7:0]) +
	( 11'sd 801) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10405) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31664) * $signed(input_fmap_77[7:0]) +
	( 14'sd 8035) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12399) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12682) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20586) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10710) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3870) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16140) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5108) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6083) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18782) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24261) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23357) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7924) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30934) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_93[7:0]) +
	( 10'sd 274) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2916) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8786) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31742) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12101) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29213) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29308) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22342) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19234) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12842) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31788) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4451) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21455) * $signed(input_fmap_113[7:0]) +
	( 11'sd 887) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10391) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19124) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19648) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17997) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13788) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 15'sd 8554) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19550) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17065) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27826) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9204) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2762) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6658) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26805) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21774) * $signed(input_fmap_13[7:0]) +
	( 10'sd 387) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31152) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15845) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16927) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31811) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11937) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11505) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13091) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9814) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18614) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26940) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14870) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23087) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13225) * $signed(input_fmap_36[7:0]) +
	( 11'sd 770) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8173) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31177) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6093) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18788) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7773) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6696) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23651) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31215) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21849) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26511) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1194) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12756) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31682) * $signed(input_fmap_56[7:0]) +
	( 11'sd 575) * $signed(input_fmap_57[7:0]) +
	( 8'sd 98) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22948) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22129) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7610) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20851) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20171) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24004) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9915) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20357) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9795) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3514) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25153) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31245) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3773) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19219) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2355) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22758) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11782) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22439) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16921) * $signed(input_fmap_97[7:0]) +
	( 12'sd 2023) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23002) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15311) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25854) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9901) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1390) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18793) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4401) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29336) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3420) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8728) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23088) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1997) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7838) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26576) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3826) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9190) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24574) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19438) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11812) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26845) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19560) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 16'sd 22244) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16392) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24669) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10218) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10310) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10664) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9001) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8621) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32482) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15974) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1331) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4323) * $signed(input_fmap_20[7:0]) +
	( 5'sd 13) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30536) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14380) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6738) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4981) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14237) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28509) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22536) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25303) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23000) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11865) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18659) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30393) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11708) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18115) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8842) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30508) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20808) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29833) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6514) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14106) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2912) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25493) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21306) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20272) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13090) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2170) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28322) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9818) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29674) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21378) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23826) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5686) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5560) * $signed(input_fmap_65[7:0]) +
	( 11'sd 929) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31085) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4528) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26852) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9353) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13123) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12829) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24494) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13323) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24636) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3060) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12483) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_88[7:0]) +
	( 11'sd 744) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10497) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10032) * $signed(input_fmap_95[7:0]) +
	( 14'sd 8115) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31355) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21339) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29110) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13358) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2344) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12375) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4240) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25342) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30749) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32348) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28401) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6964) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14066) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18440) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17669) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19721) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24163) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32716) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21867) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7747) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14858) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 16'sd 26597) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7816) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6122) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11839) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21911) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7878) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9772) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23854) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29186) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32417) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17629) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13987) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13836) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13449) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22906) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2580) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18901) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13975) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4722) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18173) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14516) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5751) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19937) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30849) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21515) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23542) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24029) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19783) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17863) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13929) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12695) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13035) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24978) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31105) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5754) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21886) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23570) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29908) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13269) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24097) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22317) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12820) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1387) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2894) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30844) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_83[7:0]) +
	( 9'sd 157) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11246) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13861) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14763) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10859) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11545) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17299) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31956) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_102[7:0]) +
	( 11'sd 912) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23600) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26450) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20267) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14128) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6282) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14931) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17540) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31331) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12329) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_115[7:0]) +
	( 10'sd 487) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18385) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30936) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29480) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20068) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11563) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 16'sd 18488) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32345) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21665) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13159) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29292) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8918) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17591) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7150) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6174) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19491) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15293) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5079) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18869) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22153) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3492) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21844) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1740) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3147) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25230) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6714) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6933) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29057) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7775) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20022) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2088) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14860) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26306) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30457) * $signed(input_fmap_37[7:0]) +
	( 13'sd 4079) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10010) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2965) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19107) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19508) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28365) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3356) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12845) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14716) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5138) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13784) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1544) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19198) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15826) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26769) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13239) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32299) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25775) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3314) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14814) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6353) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16977) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6372) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30873) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16212) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6691) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12079) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5945) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1341) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8930) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26248) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7370) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32456) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16962) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_84[7:0]) +
	( 11'sd 968) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15690) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11598) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29286) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1710) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23195) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15413) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11555) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2968) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26947) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9683) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26524) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24909) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22614) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31396) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27716) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27812) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5285) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_115[7:0]) +
	( 10'sd 337) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29809) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13592) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5962) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6097) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15913) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6154) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24066) * $signed(input_fmap_124[7:0]) +
	( 10'sd 479) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32073) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29403) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 13'sd 3960) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14867) * $signed(input_fmap_1[7:0]) +
	( 11'sd 864) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17653) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31020) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17023) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20558) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4969) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32747) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29549) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7139) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4126) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16560) * $signed(input_fmap_15[7:0]) +
	( 12'sd 2018) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19015) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10374) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3908) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31412) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9615) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21506) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26840) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8366) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18310) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18230) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32444) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3313) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16616) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13054) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13409) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26464) * $signed(input_fmap_43[7:0]) +
	( 10'sd 326) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11892) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_48[7:0]) +
	( 11'sd 965) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17597) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2525) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26786) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30340) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21411) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31005) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25493) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11084) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17458) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19739) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15600) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23147) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3227) * $signed(input_fmap_73[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28114) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30859) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24213) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7762) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18256) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8491) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13080) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16029) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24271) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14358) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11664) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9238) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_97[7:0]) +
	( 10'sd 495) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18562) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24839) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4450) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23312) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31115) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3725) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6816) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9987) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25938) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15851) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24275) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6116) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31479) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 15'sd 12696) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6050) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1396) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27144) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14474) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16253) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27545) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21235) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6074) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1338) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4230) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4421) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14967) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22185) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28867) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7215) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8219) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8138) * $signed(input_fmap_29[7:0]) +
	( 10'sd 438) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19415) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31347) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10164) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14836) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28526) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13751) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5960) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16406) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14859) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29135) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16334) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31860) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21442) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12621) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28954) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10931) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22363) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17628) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13782) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23948) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13827) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27542) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28658) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31465) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11856) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1659) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5558) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21451) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20838) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10381) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13044) * $signed(input_fmap_80[7:0]) +
	( 10'sd 356) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8279) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31479) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12826) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5255) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5362) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28051) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12757) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8315) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30404) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9624) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20599) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6649) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2598) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3349) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16218) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5922) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2465) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3190) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28089) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24045) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5443) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11708) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30339) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8605) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16754) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28405) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18213) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28518) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6405) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 13'sd 4077) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31302) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2365) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16474) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17005) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14635) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17224) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15319) * $signed(input_fmap_11[7:0]) +
	( 11'sd 984) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4820) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28391) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16813) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12229) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23294) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16542) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20043) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10719) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4563) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22979) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17891) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1884) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19739) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20084) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29633) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8618) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31660) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8676) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28138) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13457) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12547) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21923) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8803) * $signed(input_fmap_50[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20011) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12582) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16067) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19991) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22320) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5921) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19768) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27220) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9896) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6244) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15270) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22037) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14186) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31853) * $signed(input_fmap_77[7:0]) +
	( 11'sd 591) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19095) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1466) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5905) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3721) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2235) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9770) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15430) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1316) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_89[7:0]) +
	( 10'sd 376) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29561) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13305) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26430) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14838) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22558) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11645) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31531) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32586) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24453) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20940) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20116) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7598) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27416) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7622) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12087) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4687) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11489) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4175) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2582) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27869) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11173) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 10'sd 278) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28125) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14260) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22377) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20747) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13411) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1308) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4679) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27852) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6346) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22450) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5586) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21027) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5645) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22209) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26247) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15352) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4374) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25163) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19537) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7434) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18565) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5775) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7001) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17360) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21912) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17800) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30079) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22240) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5497) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11084) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13740) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28555) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2569) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6937) * $signed(input_fmap_54[7:0]) +
	( 10'sd 481) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10052) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4979) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17923) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21949) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23626) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18346) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16932) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30735) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28209) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1610) * $signed(input_fmap_67[7:0]) +
	( 11'sd 756) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24822) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_71[7:0]) +
	( 10'sd 326) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28091) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20542) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30362) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9465) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25818) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_79[7:0]) +
	( 8'sd 88) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15709) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26053) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32717) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26336) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19468) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21962) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23297) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2836) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25111) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6284) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25935) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19070) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29718) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13638) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6344) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20022) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_99[7:0]) +
	( 9'sd 255) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6903) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13330) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13551) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14150) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2960) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10922) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19345) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20855) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10946) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6388) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29738) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26326) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1720) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 15'sd 11089) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22466) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10706) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21622) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8825) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25272) * $signed(input_fmap_8[7:0]) +
	( 11'sd 727) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30827) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12372) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27304) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4114) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25547) * $signed(input_fmap_17[7:0]) +
	( 10'sd 457) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10453) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27371) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3265) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23574) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21199) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25710) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22493) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26532) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3843) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5334) * $signed(input_fmap_32[7:0]) +
	( 9'sd 195) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3306) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18726) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23109) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17189) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2689) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13434) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26238) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4580) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25985) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20562) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9297) * $signed(input_fmap_50[7:0]) +
	( 10'sd 404) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1512) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6801) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26838) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25800) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22788) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9630) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5158) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8799) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13006) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11885) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2756) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3921) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13375) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30947) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6421) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_77[7:0]) +
	( 7'sd 33) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2950) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12882) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18214) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5353) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3681) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16743) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18401) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25534) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_98[7:0]) +
	( 11'sd 546) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25912) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14657) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7344) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15693) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5741) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15774) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13081) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6705) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1698) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16782) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19017) * $signed(input_fmap_117[7:0]) +
	( 4'sd 6) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29634) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11520) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10129) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21977) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11078) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23672) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 14'sd 4999) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14731) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12613) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12341) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15088) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2364) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30796) * $signed(input_fmap_10[7:0]) +
	( 7'sd 53) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_12[7:0]) +
	( 11'sd 794) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24160) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4502) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3076) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20285) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11701) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18468) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5689) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30362) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2107) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16182) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9808) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16036) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19094) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26143) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32632) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22898) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_36[7:0]) +
	( 11'sd 668) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_38[7:0]) +
	( 10'sd 466) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_41[7:0]) +
	( 10'sd 274) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21671) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_44[7:0]) +
	( 11'sd 603) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24018) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9074) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21823) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10530) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29520) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10693) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21165) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6840) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31149) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22602) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5005) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28096) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19550) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12555) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22806) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_68[7:0]) +
	( 11'sd 565) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30218) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21486) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27206) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16467) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_78[7:0]) +
	( 6'sd 21) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10418) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9013) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22255) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12192) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19023) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1218) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1479) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21204) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18040) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11927) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26933) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13785) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26902) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9895) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17247) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20827) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23665) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29364) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5824) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12934) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17500) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5137) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4200) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12525) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24847) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12143) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16677) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28931) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7530) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9152) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23853) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9494) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22983) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 14'sd 6442) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8812) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_3[7:0]) +
	( 10'sd 352) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32466) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10012) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14271) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24022) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24955) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23088) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11931) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16324) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16250) * $signed(input_fmap_18[7:0]) +
	( 11'sd 620) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28773) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4574) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6054) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18530) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13290) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1051) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17270) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31806) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6911) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3646) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7878) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16856) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25084) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27312) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19065) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1516) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4482) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15185) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26307) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10347) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25175) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8888) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3470) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25822) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15135) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21628) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12134) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9891) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1864) * $signed(input_fmap_82[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25624) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11921) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11766) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16098) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18292) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31014) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13349) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23644) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14021) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7660) * $signed(input_fmap_98[7:0]) +
	( 13'sd 4027) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_101[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25704) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31530) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14182) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_110[7:0]) +
	( 15'sd 16278) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19000) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31708) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4733) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22334) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11025) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18031) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29788) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7799) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21420) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15259) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17505) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 16'sd 19351) * $signed(input_fmap_0[7:0]) +
	( 11'sd 967) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6210) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10553) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3195) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14882) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12106) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16441) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19441) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28727) * $signed(input_fmap_12[7:0]) +
	( 11'sd 593) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21917) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12635) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23134) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18725) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27739) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11215) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20323) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9711) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28223) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7576) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14307) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20186) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22718) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21326) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22719) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7319) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10336) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18154) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3468) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7027) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4569) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9124) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18071) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31005) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22095) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18200) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7633) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26826) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19569) * $signed(input_fmap_54[7:0]) +
	( 10'sd 295) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4276) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7390) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4279) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1295) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9980) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31918) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_66[7:0]) +
	( 10'sd 463) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12236) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19283) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15205) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3461) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15309) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3379) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21414) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7386) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1988) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15158) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17411) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6857) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9828) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13904) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9274) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28142) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18238) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10995) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22784) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1613) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26082) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11725) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23215) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7535) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17029) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9274) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14674) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31947) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32389) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6698) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10053) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23502) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5508) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18686) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31497) * $signed(input_fmap_121[7:0]) +
	( 8'sd 87) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31574) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 16'sd 23050) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22979) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2284) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16990) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9771) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16826) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31859) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17971) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18052) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14744) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9550) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12794) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21616) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9917) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7295) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5739) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21602) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24192) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21274) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31023) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6719) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9452) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6039) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3705) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_37[7:0]) +
	( 13'sd 4003) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16935) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13778) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30221) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31661) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6594) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22751) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22242) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28774) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20476) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5945) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19798) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15429) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25646) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14581) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18820) * $signed(input_fmap_57[7:0]) +
	( 14'sd 8129) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31364) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28279) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28718) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26179) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21127) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10941) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20257) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29188) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31549) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8815) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9811) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22435) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31731) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5032) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4871) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17852) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16122) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10560) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18432) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11386) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6667) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10737) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22841) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5518) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32340) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12763) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9042) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20316) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30086) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28489) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17129) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28910) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9732) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5795) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2500) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8319) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16273) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32349) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_121[7:0]) +
	( 10'sd 441) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16891) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20463) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 13'sd 4003) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29539) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4385) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31178) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2815) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4629) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10351) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27774) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23090) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22058) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2699) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6750) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29538) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14026) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12864) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5697) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13652) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17637) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6233) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27281) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9602) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31244) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11273) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31536) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22863) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6316) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23821) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28927) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6472) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17963) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26626) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26810) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30528) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26318) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7399) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28552) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18048) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30882) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29505) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30594) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19930) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5639) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5764) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9333) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9077) * $signed(input_fmap_64[7:0]) +
	( 9'sd 129) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22241) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31902) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9996) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10339) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25157) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5676) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7525) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9132) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7432) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29034) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31521) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6429) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12549) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9445) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21451) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6844) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10707) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29960) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17416) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21478) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16307) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_103[7:0]) +
	( 9'sd 131) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18064) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30151) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16561) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30512) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9095) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24652) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17722) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11877) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28002) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28501) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1412) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31710) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19888) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 16'sd 22164) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10528) * $signed(input_fmap_1[7:0]) +
	( 13'sd 4069) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30635) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14616) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8650) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30317) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1554) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5593) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23372) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28804) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3077) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32198) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8186) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21742) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18282) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7078) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2434) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6537) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1261) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31522) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22902) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25366) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32185) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13471) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19207) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_42[7:0]) +
	( 10'sd 484) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7399) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7820) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5153) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3809) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8486) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31802) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4554) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6954) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3003) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11055) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5891) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28292) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26790) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11308) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16292) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26822) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31153) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2285) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25390) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31304) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8291) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32010) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2862) * $signed(input_fmap_84[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10039) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23985) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7742) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_92[7:0]) +
	( 11'sd 899) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_99[7:0]) +
	( 13'sd 4070) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13528) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28213) * $signed(input_fmap_102[7:0]) +
	( 10'sd 333) * $signed(input_fmap_103[7:0]) +
	( 14'sd 8148) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24144) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12836) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9676) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5590) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7859) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24509) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7700) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9522) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2269) * $signed(input_fmap_116[7:0]) +
	( 10'sd 377) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13039) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24635) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9304) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19573) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 15'sd 13484) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16467) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11863) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24757) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13592) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12859) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23697) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30599) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20250) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32527) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25027) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16342) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6158) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5319) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2413) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25876) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24027) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24735) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6495) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2707) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10626) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24555) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26669) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29335) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28132) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9864) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16122) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4373) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16439) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13644) * $signed(input_fmap_41[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_42[7:0]) +
	( 9'sd 157) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24697) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11962) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28779) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4760) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1424) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10948) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18983) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16790) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14505) * $signed(input_fmap_57[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21143) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19411) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9809) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26385) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17044) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5085) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31840) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16282) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20798) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19029) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21152) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11609) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25267) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30473) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16883) * $signed(input_fmap_85[7:0]) +
	( 10'sd 360) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10892) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14383) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4940) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9960) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28732) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13782) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3879) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28904) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4829) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4473) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15418) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6526) * $signed(input_fmap_99[7:0]) +
	( 10'sd 466) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27090) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12474) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16756) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9128) * $signed(input_fmap_105[7:0]) +
	( 11'sd 841) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24728) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3498) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10647) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3555) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25173) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5357) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13168) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31167) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27760) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29274) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_128;
assign conv_mac_128 = 
	( 16'sd 18920) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9857) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18874) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14655) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27615) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12144) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19241) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2827) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27608) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29480) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7155) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26735) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15731) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8886) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26331) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3096) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4740) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1139) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3614) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10066) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8237) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28783) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9531) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7342) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26026) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_37[7:0]) +
	( 10'sd 473) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9779) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27897) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22420) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4150) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21533) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14441) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12590) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32762) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26732) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12695) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32534) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32114) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11570) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14496) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17253) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10031) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9518) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17452) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13503) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4667) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32575) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3790) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27250) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9973) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12028) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17971) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23876) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2381) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26046) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30350) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7207) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15574) * $signed(input_fmap_88[7:0]) +
	( 11'sd 999) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8587) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5782) * $signed(input_fmap_91[7:0]) +
	( 10'sd 416) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14918) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13306) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3958) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20473) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1414) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29623) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2437) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10448) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11807) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18994) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7439) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30183) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9083) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28856) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6752) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16019) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32049) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7827) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21890) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12009) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31279) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_129;
assign conv_mac_129 = 
	( 16'sd 30021) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3293) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2752) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13515) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22832) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31777) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3522) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11762) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24452) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24642) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21675) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18992) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7501) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6093) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3557) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15509) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21596) * $signed(input_fmap_25[7:0]) +
	( 11'sd 997) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5774) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7856) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9316) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5275) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9289) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31133) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20900) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32747) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3020) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2321) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2266) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21035) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6230) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27903) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4171) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6754) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15096) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14697) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32057) * $signed(input_fmap_63[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13109) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25116) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_69[7:0]) +
	( 11'sd 861) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26901) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15948) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21416) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26943) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16567) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29982) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31919) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31094) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1809) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22657) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18125) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17466) * $signed(input_fmap_90[7:0]) +
	( 14'sd 8059) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31509) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1189) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10545) * $signed(input_fmap_95[7:0]) +
	( 11'sd 1016) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7807) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16058) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5762) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30150) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6009) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31997) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32499) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21146) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13224) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21008) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23783) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10788) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30352) * $signed(input_fmap_114[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3913) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24753) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3262) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9164) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19705) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27068) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_130;
assign conv_mac_130 = 
	( 16'sd 23295) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27020) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8273) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28724) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20505) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19374) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9753) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15400) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20666) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10898) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22226) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_22[7:0]) +
	( 10'sd 489) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28705) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27210) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30885) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20979) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7884) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25613) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8676) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24442) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15262) * $signed(input_fmap_39[7:0]) +
	( 11'sd 955) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7859) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19326) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11505) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14744) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_45[7:0]) +
	( 11'sd 670) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26835) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25581) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3516) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11250) * $signed(input_fmap_50[7:0]) +
	( 11'sd 980) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1181) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30506) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14494) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22028) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26083) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1471) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13020) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19333) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31583) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26406) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9038) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18659) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18694) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17835) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9913) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16201) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23832) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19318) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11087) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_81[7:0]) +
	( 10'sd 460) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_85[7:0]) +
	( 14'sd 8012) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6496) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19086) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24277) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4100) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24250) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10989) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12381) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13735) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32671) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15069) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29927) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7304) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26475) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22171) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16719) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10069) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13862) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3601) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22990) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12296) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9700) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4272) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9316) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_125[7:0]) +
	( 9'sd 156) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1343) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_131;
assign conv_mac_131 = 
	( 16'sd 19014) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30865) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27655) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21100) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8897) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14968) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7821) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12577) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21747) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2458) * $signed(input_fmap_13[7:0]) +
	( 10'sd 364) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29005) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16277) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8875) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4851) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25537) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1796) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26749) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11846) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6538) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10017) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4794) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20843) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17338) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2309) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22617) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15937) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2536) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9159) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7247) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_45[7:0]) +
	( 10'sd 406) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19670) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30749) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29827) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24158) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_55[7:0]) +
	( 8'sd 125) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21843) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10170) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8010) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30831) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16925) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13465) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32148) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18354) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26496) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27946) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17063) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12130) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32419) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23295) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6962) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11384) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11212) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17151) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11992) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22469) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19736) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29257) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18035) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17550) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3144) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14513) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26329) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10770) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7936) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_101[7:0]) +
	( 11'sd 790) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25280) * $signed(input_fmap_103[7:0]) +
	( 10'sd 310) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17124) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10387) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23633) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24598) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5814) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31264) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25295) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24463) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19220) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2630) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2123) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24270) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22581) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_122[7:0]) +
	( 11'sd 767) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27022) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25093) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_132;
assign conv_mac_132 = 
	( 15'sd 8345) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3012) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12005) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1679) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_4[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23417) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29883) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5142) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18498) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19490) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32175) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28197) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16546) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11628) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5872) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1056) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17634) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25355) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13086) * $signed(input_fmap_26[7:0]) +
	( 11'sd 825) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19495) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7691) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27099) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1890) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12421) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8680) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3767) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2774) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6406) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8549) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28102) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21528) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23906) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21399) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12980) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17447) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22768) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6283) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23934) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9543) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12895) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16786) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22871) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10313) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13198) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1997) * $signed(input_fmap_66[7:0]) +
	( 13'sd 4030) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6521) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23599) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3585) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11233) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22339) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21045) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29539) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17412) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5988) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8698) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20578) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14812) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28992) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_85[7:0]) +
	( 11'sd 933) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3620) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16874) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11556) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1736) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8996) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6526) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32482) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28838) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21931) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29246) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32520) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18424) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10946) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24521) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10293) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18338) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17873) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18641) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11959) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15635) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18089) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3351) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_133;
assign conv_mac_133 = 
	( 16'sd 22918) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31627) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27982) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26412) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1214) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21077) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22754) * $signed(input_fmap_6[7:0]) +
	( 10'sd 360) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22649) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18511) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15208) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22463) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30008) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7197) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5795) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24853) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21766) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8084) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14826) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16547) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13982) * $signed(input_fmap_28[7:0]) +
	( 11'sd 630) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30153) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20422) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26216) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2559) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25761) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27350) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16211) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7941) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27231) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1572) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10024) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22650) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20339) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2761) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9091) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4926) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13949) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27099) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15243) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15068) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24955) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27209) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20412) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31239) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27789) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13334) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18074) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8956) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8534) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4511) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23487) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25455) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32629) * $signed(input_fmap_80[7:0]) +
	( 11'sd 541) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23054) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8272) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13987) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8923) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7688) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3553) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15814) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12675) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31286) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31373) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3675) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32701) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14928) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14473) * $signed(input_fmap_107[7:0]) +
	( 10'sd 341) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18297) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13865) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13099) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9003) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14251) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29746) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6590) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19610) * $signed(input_fmap_118[7:0]) +
	( 10'sd 363) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16447) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29310) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14212) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32622) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14054) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11101) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_134;
assign conv_mac_134 = 
	( 16'sd 28195) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19902) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4399) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14370) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8946) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5297) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8956) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2887) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23822) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9125) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27977) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12899) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23123) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17775) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20623) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20527) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14070) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26027) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13812) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23294) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31511) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28322) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11885) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30811) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14770) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17388) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31170) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5337) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1908) * $signed(input_fmap_45[7:0]) +
	( 9'sd 255) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29530) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31675) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19223) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10004) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8734) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21991) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7546) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29107) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6475) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29236) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7369) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4119) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14725) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22755) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12545) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7485) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8959) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14955) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22393) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24873) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28743) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20221) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17907) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20019) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_83[7:0]) +
	( 11'sd 926) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_87[7:0]) +
	( 11'sd 826) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7312) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8131) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2670) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6105) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8928) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24980) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6413) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5290) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12794) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12719) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29943) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9294) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24627) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15403) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22322) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8203) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29438) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31047) * $signed(input_fmap_118[7:0]) +
	( 11'sd 675) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17990) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10237) * $signed(input_fmap_121[7:0]) +
	( 10'sd 355) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18976) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15897) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_135;
assign conv_mac_135 = 
	( 15'sd 9560) * $signed(input_fmap_0[7:0]) +
	( 11'sd 763) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5219) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19648) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9445) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22986) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2094) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7270) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12410) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25947) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8899) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19305) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17314) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3221) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16170) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6470) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32590) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5901) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14460) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27804) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12670) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4572) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32628) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31829) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22835) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6240) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30365) * $signed(input_fmap_38[7:0]) +
	( 10'sd 312) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2855) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17910) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23331) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4643) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12825) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10338) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16436) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23978) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29310) * $signed(input_fmap_55[7:0]) +
	( 11'sd 787) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6775) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24375) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13173) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32583) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12263) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12092) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25031) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5868) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17647) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13304) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4355) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27213) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4615) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17805) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2244) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18849) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13326) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27434) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11603) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27992) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17357) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18891) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14246) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3595) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24321) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1638) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1358) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15500) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10457) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21473) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23791) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2508) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20810) * $signed(input_fmap_105[7:0]) +
	( 11'sd 940) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20186) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21870) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3796) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29515) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25354) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25809) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28974) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6239) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7730) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13944) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9294) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7498) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12892) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6417) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14610) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_136;
assign conv_mac_136 = 
	( 15'sd 13234) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16072) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15361) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18683) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15745) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16273) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20151) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25636) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21396) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1463) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19942) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24297) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23953) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20099) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4668) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4857) * $signed(input_fmap_25[7:0]) +
	( 11'sd 760) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28460) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1490) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3550) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6556) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22906) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25806) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21924) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26742) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7495) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5144) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19254) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22691) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24232) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9358) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13602) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30867) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1931) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5460) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2731) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21950) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11015) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23912) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_56[7:0]) +
	( 10'sd 276) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11109) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32467) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25888) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23071) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31243) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10298) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28072) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8810) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26243) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14931) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18935) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17152) * $signed(input_fmap_73[7:0]) +
	( 10'sd 357) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7022) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16284) * $signed(input_fmap_77[7:0]) +
	( 11'sd 727) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23282) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19263) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29909) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12486) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15170) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9667) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28277) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24547) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12059) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32526) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18868) * $signed(input_fmap_93[7:0]) +
	( 13'sd 4076) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26206) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17501) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2412) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3532) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2489) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6217) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30041) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16268) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2739) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16297) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24585) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26722) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32209) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20748) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29560) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8749) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3217) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8935) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10597) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19361) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30846) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_137;
assign conv_mac_137 = 
	( 16'sd 20654) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28575) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20259) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20625) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1797) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28001) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20107) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18685) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29717) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6844) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18208) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9009) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3210) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2324) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29978) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8615) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22028) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21395) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2405) * $signed(input_fmap_34[7:0]) +
	( 10'sd 339) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8093) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22190) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15811) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29165) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19655) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20359) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30456) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11244) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31539) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32371) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7445) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24840) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11678) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5935) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15447) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14408) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30218) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7412) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18216) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19243) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31274) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8682) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12565) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7387) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5692) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24967) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29561) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24831) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30325) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7983) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27970) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11738) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29331) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22863) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29277) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8896) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23885) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9799) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22547) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11021) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30150) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11042) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9353) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8250) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5113) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_113[7:0]) +
	( 11'sd 633) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26856) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6401) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17580) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16500) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31725) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22142) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31905) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_138;
assign conv_mac_138 = 
	( 16'sd 23176) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21432) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18717) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28777) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11664) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31700) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7582) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23673) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10117) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3323) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25127) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3787) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14333) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20205) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_18[7:0]) +
	( 11'sd 592) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_20[7:0]) +
	( 11'sd 588) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21826) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5590) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1645) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26426) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28256) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16743) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17872) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11697) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11935) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28603) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14994) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1876) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28713) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16624) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10356) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23175) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32297) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26539) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5521) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23936) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27132) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11072) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_55[7:0]) +
	( 11'sd 793) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5812) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7002) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10000) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5581) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11189) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10879) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8527) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28687) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21848) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9171) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9995) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2642) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25707) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18347) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21474) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22266) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10943) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24978) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14783) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2339) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24232) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26139) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9145) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8068) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29994) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1064) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26539) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6032) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7333) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24444) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25540) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27989) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17408) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29329) * $signed(input_fmap_115[7:0]) +
	( 11'sd 964) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29693) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18586) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3212) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18723) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30561) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_139;
assign conv_mac_139 = 
	( 12'sd 1315) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25370) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9781) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5280) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9381) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_5[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13745) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12954) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21493) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12809) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23435) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28514) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1104) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21159) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6892) * $signed(input_fmap_18[7:0]) +
	( 10'sd 496) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3516) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_22[7:0]) +
	( 13'sd 4072) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7096) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28567) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6964) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18683) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26891) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11976) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12756) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18000) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2442) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29349) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11762) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1806) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11928) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4682) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20908) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18603) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8516) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13583) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10735) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17258) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19245) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30065) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4144) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24204) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14485) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8397) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31704) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21029) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29760) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9389) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11660) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27098) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2831) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30274) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6052) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32387) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23833) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29612) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6760) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24851) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24307) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_96[7:0]) +
	( 12'sd 2012) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2614) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6585) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21671) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25136) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14253) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12687) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13576) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7922) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17352) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19962) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18185) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29231) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11834) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27751) * $signed(input_fmap_115[7:0]) +
	( 11'sd 602) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30609) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13235) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10989) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22451) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7991) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29370) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28921) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_140;
assign conv_mac_140 = 
	( 13'sd 3566) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23475) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11633) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31762) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1815) * $signed(input_fmap_7[7:0]) +
	( 9'sd 229) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23739) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16450) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31368) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25414) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27506) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21289) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25173) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6180) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_18[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9484) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22725) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29571) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19690) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5331) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3446) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3225) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7311) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11984) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6705) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25803) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30539) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3382) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25231) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3612) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13815) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11869) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10373) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22602) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29762) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15774) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23781) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19994) * $signed(input_fmap_57[7:0]) +
	( 10'sd 382) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_59[7:0]) +
	( 10'sd 332) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29309) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2620) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9436) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6044) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3217) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30229) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25079) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18423) * $signed(input_fmap_72[7:0]) +
	( 11'sd 525) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4184) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18479) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5158) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_78[7:0]) +
	( 11'sd 822) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8429) * $signed(input_fmap_80[7:0]) +
	( 13'sd 4063) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28789) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13954) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31208) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2095) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5084) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23062) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7359) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11923) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29030) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18502) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24007) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12316) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9675) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4827) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8425) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12873) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8451) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26868) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20552) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9433) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_111[7:0]) +
	( 6'sd 22) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13158) * $signed(input_fmap_113[7:0]) +
	( 13'sd 4033) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11846) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31598) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13952) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14087) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21978) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23278) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21312) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23035) * $signed(input_fmap_124[7:0]) +
	( 11'sd 895) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_126[7:0]) +
	( 10'sd 391) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_141;
assign conv_mac_141 = 
	( 15'sd 13457) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10437) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8978) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5762) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20461) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31548) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19669) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14329) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4986) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29333) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12798) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6467) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15722) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20235) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3753) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28430) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28717) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10437) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14881) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21399) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30943) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19904) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12775) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10780) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16814) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20148) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9730) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26186) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29814) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32638) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17723) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2280) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4483) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27834) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3432) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29978) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29027) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20420) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_63[7:0]) +
	( 17'sd 32768) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10894) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27037) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12303) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11483) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26253) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22761) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11508) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8934) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13286) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23092) * $signed(input_fmap_77[7:0]) +
	( 14'sd 8075) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7944) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31024) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14141) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8543) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17547) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15585) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20149) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23311) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4692) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22728) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27431) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15500) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5623) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8798) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16605) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19836) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22298) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9173) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9104) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23699) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30657) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7410) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_142;
assign conv_mac_142 = 
	( 13'sd 3392) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_1[7:0]) +
	( 13'sd 4007) * $signed(input_fmap_2[7:0]) +
	( 11'sd 676) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29416) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1805) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26796) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1913) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26394) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11226) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14487) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9746) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10588) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24357) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8660) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12553) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19945) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30881) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28232) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3070) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5789) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15560) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18276) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30412) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7804) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31298) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24853) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7816) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17135) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30649) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8907) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9883) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3431) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5253) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2985) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18984) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12121) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31246) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23469) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30798) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11397) * $signed(input_fmap_64[7:0]) +
	( 11'sd 569) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12827) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7500) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3783) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29487) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9366) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21695) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10715) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8408) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14255) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13703) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11609) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31014) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2427) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11448) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20909) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23459) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15255) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31593) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14169) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3767) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21939) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_95[7:0]) +
	( 11'sd 660) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22005) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1030) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29113) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21724) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3455) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14257) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21436) * $signed(input_fmap_103[7:0]) +
	( 11'sd 751) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17173) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7180) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31041) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26864) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14080) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5204) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14155) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12526) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9659) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18580) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1122) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4385) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27784) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14563) * $signed(input_fmap_125[7:0]) +
	( 15'sd 16369) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_143;
assign conv_mac_143 = 
	( 16'sd 20557) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6330) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_2[7:0]) +
	( 11'sd 908) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16412) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32649) * $signed(input_fmap_8[7:0]) +
	( 11'sd 762) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31471) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11363) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24286) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20977) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15910) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14313) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19801) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14611) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_27[7:0]) +
	( 11'sd 515) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11006) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18702) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5093) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20802) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5154) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19105) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32425) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11569) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1033) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14132) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_42[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28368) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9039) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5014) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7850) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25455) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22335) * $signed(input_fmap_50[7:0]) +
	( 11'sd 868) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11205) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15075) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11334) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31463) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23487) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1035) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31274) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20073) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25477) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6600) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_65[7:0]) +
	( 11'sd 686) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10209) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2827) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22270) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6671) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24911) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24184) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14666) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17686) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2778) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16608) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28549) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24853) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14596) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8511) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16604) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13482) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20954) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18754) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18289) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_98[7:0]) +
	( 10'sd 272) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7640) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9324) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14481) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30527) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11925) * $signed(input_fmap_107[7:0]) +
	( 11'sd 669) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4700) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3408) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31561) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11988) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9377) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31618) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6396) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28875) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_144;
assign conv_mac_144 = 
	( 16'sd 19777) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3125) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25285) * $signed(input_fmap_2[7:0]) +
	( 11'sd 729) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4192) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18493) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1547) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18852) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20247) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22031) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20486) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11619) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14392) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11934) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3741) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28103) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17960) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2813) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4860) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13025) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22897) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30376) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5380) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31552) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17323) * $signed(input_fmap_30[7:0]) +
	( 14'sd 8102) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3710) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1219) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29620) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9155) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15326) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28057) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11457) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15664) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22871) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29016) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16723) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9504) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31443) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16684) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29255) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26211) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29056) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30464) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30694) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14055) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28476) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32283) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17314) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1035) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1587) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12156) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13802) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25154) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10487) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28793) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10033) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7105) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26974) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16968) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30311) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18267) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19121) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29080) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2715) * $signed(input_fmap_92[7:0]) +
	( 8'sd 68) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14691) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29172) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12121) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16317) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3748) * $signed(input_fmap_100[7:0]) +
	( 11'sd 882) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6174) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9527) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11440) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7895) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4774) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30572) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22091) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_115[7:0]) +
	( 10'sd 288) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_118[7:0]) +
	( 6'sd 30) * $signed(input_fmap_119[7:0]) +
	( 11'sd 536) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13309) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4409) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24840) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30155) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7727) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_145;
assign conv_mac_145 = 
	( 16'sd 22430) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31119) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28498) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3505) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14298) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11478) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4287) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13618) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4648) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10264) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_15[7:0]) +
	( 10'sd 319) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7919) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20045) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19323) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8147) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13825) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8344) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8282) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18861) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23891) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17314) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26709) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2532) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15393) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26228) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10241) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31410) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13501) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21153) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5558) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5419) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30995) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2331) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32557) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13774) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16244) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11203) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13713) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_66[7:0]) +
	( 11'sd 529) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20447) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4468) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21894) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17426) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16246) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25019) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10215) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9702) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16615) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11529) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5560) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2413) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13833) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9273) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26158) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4726) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18852) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2101) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18917) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11830) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22130) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_110[7:0]) +
	( 9'sd 141) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9921) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23817) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10782) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13842) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28388) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18747) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30103) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13848) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14585) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8112) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_146;
assign conv_mac_146 = 
	( 13'sd 2237) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23359) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2632) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9841) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6694) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13958) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21339) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18796) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16027) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28960) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32404) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30021) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13009) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7797) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29028) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24895) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14321) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4337) * $signed(input_fmap_29[7:0]) +
	( 11'sd 809) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2248) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25979) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13168) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14477) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20910) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5160) * $signed(input_fmap_40[7:0]) +
	( 10'sd 343) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15834) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11480) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22304) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3246) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5280) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4504) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18738) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10808) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8917) * $signed(input_fmap_50[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13848) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15050) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17318) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5960) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13644) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1641) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16520) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7666) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23043) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31802) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_73[7:0]) +
	( 11'sd 913) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32579) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1563) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26216) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17766) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3372) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31079) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30145) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11989) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4460) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17879) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27240) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26846) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1935) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26692) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11414) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1385) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17367) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12919) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4709) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8203) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24521) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21057) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10432) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12162) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7054) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12910) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31983) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18195) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5038) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6127) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14671) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7880) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19132) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20105) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30092) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10789) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_147;
assign conv_mac_147 = 
	( 16'sd 19781) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15822) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23932) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8629) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13732) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10421) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32040) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13170) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3394) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14770) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8505) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6014) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10472) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15465) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3610) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10959) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20424) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5826) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20861) * $signed(input_fmap_34[7:0]) +
	( 7'sd 41) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12410) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18347) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23976) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21216) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5743) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21579) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28763) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24346) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13841) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32597) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23237) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1286) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8040) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25845) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2460) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23880) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21086) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1175) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16874) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22371) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_72[7:0]) +
	( 11'sd 685) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19852) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13835) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19307) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10547) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15119) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24082) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13951) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26343) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_92[7:0]) +
	( 11'sd 688) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9024) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28475) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3124) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11091) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11364) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31905) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2699) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32449) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29288) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11572) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14230) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21408) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17764) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17245) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30230) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5708) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12475) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32570) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_117[7:0]) +
	( 11'sd 573) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4104) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2775) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32418) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19278) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28186) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9961) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31226) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_148;
assign conv_mac_148 = 
	( 16'sd 23013) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21015) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30130) * $signed(input_fmap_2[7:0]) +
	( 11'sd 738) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10311) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3251) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17920) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30744) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21743) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2752) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32180) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22427) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3556) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10188) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17407) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29460) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9706) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17746) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24143) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11899) * $signed(input_fmap_28[7:0]) +
	( 10'sd 337) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12900) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1618) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12787) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4096) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1093) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4421) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6367) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9461) * $signed(input_fmap_40[7:0]) +
	( 11'sd 856) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17554) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3351) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21270) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24015) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5847) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_49[7:0]) +
	( 12'sd 2002) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12593) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1352) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21404) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25861) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18597) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24810) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11703) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9195) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31572) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23925) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13262) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8610) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6142) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20207) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18794) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21202) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15775) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8316) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26751) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9579) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3167) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16733) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14495) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6447) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10108) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11239) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10850) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27405) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14054) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19904) * $signed(input_fmap_106[7:0]) +
	( 11'sd 965) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1951) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19867) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2984) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19738) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6175) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8275) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28692) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28777) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23647) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4741) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4175) * $signed(input_fmap_121[7:0]) +
	( 11'sd 769) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26007) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_149;
assign conv_mac_149 = 
	( 14'sd 4845) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16100) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16464) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18416) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25455) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1664) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2899) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1156) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8383) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25567) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24657) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21726) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15919) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20116) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29847) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28634) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30415) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20001) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7020) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2720) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6081) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11243) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15359) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7633) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22309) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9141) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29244) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_39[7:0]) +
	( 11'sd 948) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6987) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24172) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17191) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11435) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10213) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13499) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5756) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7130) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32163) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5355) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28861) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24811) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2112) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11361) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17121) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30527) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29833) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28037) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8164) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29098) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12094) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10974) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25950) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29471) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3380) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29059) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23509) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26446) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4429) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8718) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22080) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29582) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13327) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3118) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12325) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20460) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10126) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11634) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17790) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14398) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32628) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12319) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3308) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28152) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17231) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10795) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26865) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9644) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27876) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30386) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23042) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5772) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27388) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10921) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24757) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22472) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27193) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_150;
assign conv_mac_150 = 
	( 15'sd 13484) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21339) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20140) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9976) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25995) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5290) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23959) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22950) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28824) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27468) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15208) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2334) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4898) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25218) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21554) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2917) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21733) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14196) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28077) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23807) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20328) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2895) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18572) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26479) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15713) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16200) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23584) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8801) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16662) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5617) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6824) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19425) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24252) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1524) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3676) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3757) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10035) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25800) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18465) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4433) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21828) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32678) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14957) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25252) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21253) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22292) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29868) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31035) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7213) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30383) * $signed(input_fmap_81[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30932) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1178) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_86[7:0]) +
	( 6'sd 30) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20605) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14177) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20021) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7263) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24902) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19657) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_100[7:0]) +
	( 8'sd 125) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10913) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10083) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29066) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19692) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12057) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7419) * $signed(input_fmap_113[7:0]) +
	( 11'sd 794) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19036) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20285) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24397) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21546) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28414) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28796) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31881) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30956) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_151;
assign conv_mac_151 = 
	( 15'sd 16154) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21700) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16030) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18323) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3732) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14261) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7201) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23467) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29935) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13521) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14303) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7223) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31991) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26990) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6355) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11471) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8902) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2449) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26918) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21423) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17387) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28325) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_29[7:0]) +
	( 9'sd 198) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25794) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13361) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10514) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12779) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22055) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14941) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14183) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28699) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32082) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9234) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32242) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32026) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23180) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32565) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_52[7:0]) +
	( 10'sd 367) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5926) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_56[7:0]) +
	( 11'sd 856) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2791) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2305) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15375) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_63[7:0]) +
	( 11'sd 670) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1365) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19386) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13189) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12783) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26605) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32213) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23408) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3098) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7432) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8802) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3561) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12375) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29041) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26577) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24021) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23409) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8893) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_97[7:0]) +
	( 10'sd 342) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30230) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5010) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16769) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2775) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7576) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11558) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5633) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9855) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15622) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8787) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6630) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6383) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22237) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11330) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8767) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10975) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20953) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19826) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20659) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_152;
assign conv_mac_152 = 
	( 16'sd 17398) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5255) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30211) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14140) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11466) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30875) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30591) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28089) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11224) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_15[7:0]) +
	( 11'sd 787) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18582) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3595) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9493) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26200) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5313) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25018) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13466) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32084) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9448) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20893) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13663) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11360) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13551) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14011) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17724) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26094) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32371) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19903) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10548) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17116) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4325) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18687) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32003) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15857) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1930) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4451) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18557) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2509) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19421) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4267) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17194) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20032) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15027) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14839) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16895) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28361) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31052) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_71[7:0]) +
	( 11'sd 851) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11387) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8642) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28504) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6549) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21177) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20644) * $signed(input_fmap_82[7:0]) +
	( 10'sd 351) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8382) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24298) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11212) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21385) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31541) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8534) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30291) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5465) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21097) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12022) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30147) * $signed(input_fmap_99[7:0]) +
	( 11'sd 850) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1166) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10707) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5553) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29951) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3206) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10919) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31561) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2894) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19699) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9770) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9863) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7702) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27377) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12300) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29346) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22409) * $signed(input_fmap_120[7:0]) +
	( 12'sd 2046) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25720) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27383) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28636) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20845) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_153;
assign conv_mac_153 = 
	( 15'sd 14103) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3809) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18202) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_3[7:0]) +
	( 9'sd 251) * $signed(input_fmap_4[7:0]) +
	( 11'sd 951) * $signed(input_fmap_5[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7925) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22290) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10946) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3218) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4263) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30323) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27631) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4249) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17226) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25549) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14734) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2858) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26033) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14178) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26450) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18557) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28951) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5819) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18237) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16415) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19124) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21459) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9260) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15069) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30385) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27082) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16204) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12171) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_54[7:0]) +
	( 6'sd 23) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17419) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1033) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14589) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4544) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_66[7:0]) +
	( 14'sd 8077) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19235) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15342) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21240) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20210) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19710) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4690) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23194) * $signed(input_fmap_83[7:0]) +
	( 10'sd 422) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26922) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12338) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30678) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26837) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14551) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15620) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16112) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22057) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5062) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17674) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_99[7:0]) +
	( 10'sd 432) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27845) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25788) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3081) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31743) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9794) * $signed(input_fmap_108[7:0]) +
	( 11'sd 548) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29231) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21380) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9582) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30935) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22769) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2215) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6451) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2192) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21114) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15723) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5712) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_154;
assign conv_mac_154 = 
	( 16'sd 29577) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26986) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29012) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28382) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18896) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23257) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28399) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18684) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30677) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1231) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7844) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8721) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32278) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5794) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32745) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31606) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17959) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_31[7:0]) +
	( 10'sd 402) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7617) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8989) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31086) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24408) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19152) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22696) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17741) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7803) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28003) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5179) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18731) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3133) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30875) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14985) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22305) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22090) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32537) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27149) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16992) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18167) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13261) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25238) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11241) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2906) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13391) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11936) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17401) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23987) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30972) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26627) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17366) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16740) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23606) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32341) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31793) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20721) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31906) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15679) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18987) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6243) * $signed(input_fmap_98[7:0]) +
	( 11'sd 906) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10135) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2936) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30373) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17277) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22875) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10233) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13903) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29903) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10429) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24568) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26341) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10250) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28127) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2917) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28061) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23809) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21821) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_155;
assign conv_mac_155 = 
	( 14'sd 5107) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26062) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2960) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12316) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30668) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25546) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3228) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14893) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29846) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5403) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22583) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5521) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18706) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22461) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23814) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3479) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28683) * $signed(input_fmap_26[7:0]) +
	( 10'sd 476) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11492) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20918) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27402) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11568) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10876) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27678) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14258) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23051) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13096) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10018) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22618) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26033) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_47[7:0]) +
	( 9'sd 210) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7437) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23855) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1299) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29515) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28106) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24021) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2462) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28565) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24173) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27086) * $signed(input_fmap_60[7:0]) +
	( 9'sd 182) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27830) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_68[7:0]) +
	( 11'sd 1001) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12663) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6015) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12733) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10282) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13797) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20207) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16088) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23258) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15517) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20422) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13048) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20776) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26989) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8756) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19304) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12473) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10776) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30606) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14186) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15600) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8334) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30651) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14750) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31961) * $signed(input_fmap_116[7:0]) +
	( 9'sd 217) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14989) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23131) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28486) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26090) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9657) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9288) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30715) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_156;
assign conv_mac_156 = 
	( 16'sd 18023) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13404) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20865) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11719) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25887) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16712) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6986) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2858) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4977) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32668) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6367) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31466) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29261) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29095) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5836) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28041) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32005) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3340) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3516) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1926) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18382) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11218) * $signed(input_fmap_38[7:0]) +
	( 5'sd 14) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26972) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14150) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16147) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7075) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18532) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27663) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31221) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1863) * $signed(input_fmap_52[7:0]) +
	( 11'sd 648) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7753) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16590) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17550) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22696) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31159) * $signed(input_fmap_62[7:0]) +
	( 9'sd 179) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5558) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14692) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28890) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6304) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2649) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20514) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21573) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29670) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22503) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26374) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28454) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6493) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28386) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23084) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14761) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20179) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30369) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27299) * $signed(input_fmap_91[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28207) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31736) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6360) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2491) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31546) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20704) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16425) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4793) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29494) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28743) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29944) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25123) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20766) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6407) * $signed(input_fmap_113[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21618) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9045) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13964) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29846) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26651) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26430) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_157;
assign conv_mac_157 = 
	( 16'sd 20666) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9761) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24833) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4839) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16750) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30921) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30696) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1649) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25005) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4628) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6427) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23156) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27902) * $signed(input_fmap_20[7:0]) +
	( 12'sd 2034) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24328) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5346) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19041) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28641) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12059) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18245) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30109) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20420) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26242) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14459) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21973) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28385) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15357) * $signed(input_fmap_40[7:0]) +
	( 8'sd 79) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_42[7:0]) +
	( 10'sd 415) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3702) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25030) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26626) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5589) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_49[7:0]) +
	( 11'sd 686) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17154) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19717) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21567) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12515) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20962) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4283) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31552) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7489) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4780) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14008) * $signed(input_fmap_66[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26161) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5517) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28919) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15882) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3019) * $signed(input_fmap_74[7:0]) +
	( 7'sd 42) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12261) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16736) * $signed(input_fmap_78[7:0]) +
	( 10'sd 456) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29685) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2989) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17944) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16923) * $signed(input_fmap_83[7:0]) +
	( 11'sd 742) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18900) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30275) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5048) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29258) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19103) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26146) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20848) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6715) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11742) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18220) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16182) * $signed(input_fmap_100[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29748) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15313) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20623) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27978) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5132) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14784) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9296) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28706) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9922) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15202) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16065) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13489) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29508) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3282) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4512) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9013) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10082) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21099) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4810) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_158;
assign conv_mac_158 = 
	( 16'sd 32695) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14334) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20516) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14634) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24077) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23008) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13054) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5242) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14396) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9695) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9830) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9198) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32394) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18431) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20465) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28982) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30967) * $signed(input_fmap_21[7:0]) +
	( 10'sd 492) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20060) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20664) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9244) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12491) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25222) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9662) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13760) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21147) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13660) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27441) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14790) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7353) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9736) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7241) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_45[7:0]) +
	( 13'sd 4049) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3418) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21980) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2471) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17023) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9334) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22101) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11180) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8335) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11748) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6795) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11175) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24634) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30382) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30470) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14259) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15182) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24252) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5313) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32496) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32448) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29476) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31792) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9952) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10892) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26053) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14020) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_85[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10077) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6769) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2086) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19851) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22998) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6602) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2740) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31838) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26970) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3278) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16925) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6945) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19168) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6852) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7272) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2349) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13150) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5880) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29427) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16667) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19999) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14484) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13819) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19472) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_159;
assign conv_mac_159 = 
	( 16'sd 27407) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21855) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20210) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15771) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1407) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12691) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23335) * $signed(input_fmap_7[7:0]) +
	( 10'sd 324) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1728) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23676) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28789) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19875) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4803) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10144) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17716) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30485) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22239) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8524) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9495) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_24[7:0]) +
	( 8'sd 65) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14457) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2910) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_29[7:0]) +
	( 11'sd 732) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7700) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31966) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9148) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13743) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30109) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6182) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24695) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24593) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4738) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30989) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20665) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21818) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21431) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2350) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28576) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30411) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23137) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17819) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26054) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14675) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15824) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7178) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15681) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29958) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8143) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4630) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7192) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14548) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12356) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28708) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22470) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28530) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30737) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32502) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12011) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25341) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14200) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23837) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6274) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20159) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27711) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18437) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26182) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10683) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12418) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8351) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15496) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30075) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10580) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14988) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10516) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21242) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29623) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8919) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1391) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8585) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27975) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20863) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32681) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3648) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2400) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29586) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3061) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22027) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13710) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_160;
assign conv_mac_160 = 
	( 16'sd 21442) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15458) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24768) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16508) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30492) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28037) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17141) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6195) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16971) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13234) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9430) * $signed(input_fmap_17[7:0]) +
	( 8'sd 96) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10442) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13771) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21853) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7597) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24681) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3149) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1193) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19043) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17509) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7428) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7135) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31365) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9336) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1636) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29825) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29546) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5576) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23669) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12725) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24288) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23124) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9904) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18543) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28999) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_60[7:0]) +
	( 11'sd 979) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31252) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32052) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14700) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8860) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14942) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16826) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15563) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31359) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6908) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28274) * $signed(input_fmap_81[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11466) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30671) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14134) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32281) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2321) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6279) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10124) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10576) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30061) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32158) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28302) * $signed(input_fmap_101[7:0]) +
	( 8'sd 112) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_103[7:0]) +
	( 14'sd 8007) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22416) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22127) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25433) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12566) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24381) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23452) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18675) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30409) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12481) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26722) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26809) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14958) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_161;
assign conv_mac_161 = 
	( 16'sd 31138) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26103) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28576) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3713) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19682) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27269) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24999) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31774) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25313) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12495) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24384) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1781) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26731) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24850) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8183) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11480) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5369) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20217) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13928) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18309) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10716) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9427) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1878) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14757) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3872) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3454) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13609) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30900) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20089) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31423) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1676) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12407) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28977) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17956) * $signed(input_fmap_47[7:0]) +
	( 9'sd 181) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10756) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28371) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32748) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21408) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28851) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5198) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16318) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4627) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5509) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16516) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19747) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30353) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6087) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7788) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9542) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21585) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29024) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29180) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29747) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11982) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6806) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16864) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18935) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11859) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16803) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23201) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30890) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12991) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3319) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5379) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25224) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31949) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20486) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8871) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14246) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24471) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11143) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32419) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3770) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14853) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10957) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11679) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9961) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6913) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16299) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28906) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10294) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31280) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14493) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6873) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16013) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23924) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29843) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1887) * $signed(input_fmap_126[7:0]) +
	( 11'sd 544) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_162;
assign conv_mac_162 = 
	( 16'sd 18875) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13242) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16313) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10239) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16312) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26689) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7989) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29184) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22599) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19797) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9627) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28443) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27711) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8943) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8231) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14004) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30732) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7964) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19488) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3559) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12848) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32308) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7979) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24041) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25918) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15350) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27232) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27529) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23108) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8646) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9937) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31490) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7858) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15542) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19758) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15285) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19795) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30058) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14728) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27356) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4912) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1887) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21506) * $signed(input_fmap_60[7:0]) +
	( 11'sd 750) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5919) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1219) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18804) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2291) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25885) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29748) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29439) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27697) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10020) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5496) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15218) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29574) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29939) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13842) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24555) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14283) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26694) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15815) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31380) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24462) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22760) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27009) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21482) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3451) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19916) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6625) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9850) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14826) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27571) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20162) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3865) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19249) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23384) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24575) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27369) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8725) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4361) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15798) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22791) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_163;
assign conv_mac_163 = 
	( 16'sd 24640) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14106) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18225) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18529) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23656) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10455) * $signed(input_fmap_8[7:0]) +
	( 10'sd 470) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10303) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1385) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13086) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6998) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7636) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14757) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12413) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23214) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29830) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22126) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29654) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28743) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9454) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6781) * $signed(input_fmap_30[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12035) * $signed(input_fmap_32[7:0]) +
	( 9'sd 254) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5170) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29794) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13985) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7378) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15188) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32721) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2848) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30466) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_45[7:0]) +
	( 11'sd 977) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31918) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8868) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29924) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19118) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26617) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26747) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16745) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26248) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_55[7:0]) +
	( 11'sd 781) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26216) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5655) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28668) * $signed(input_fmap_61[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21712) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12080) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18173) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28488) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12823) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13622) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10057) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12754) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16637) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2266) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26957) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16802) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25104) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5266) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21780) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30561) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27416) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20610) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4839) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8804) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8461) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21378) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4162) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7210) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13956) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22795) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9666) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15084) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7157) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2553) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26779) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16834) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1408) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16164) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8491) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24913) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5142) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20597) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16240) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_125[7:0]) +
	( 14'sd 8070) * $signed(input_fmap_126[7:0]) +
	( 10'sd 381) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_164;
assign conv_mac_164 = 
	( 16'sd 31819) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31707) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12849) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29556) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22695) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22339) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2917) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18346) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28846) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31827) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30109) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2873) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7153) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12135) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15268) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5839) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18437) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32451) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9651) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15204) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5032) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29498) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23641) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24193) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13739) * $signed(input_fmap_33[7:0]) +
	( 10'sd 416) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26919) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22552) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30138) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5223) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9179) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17934) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32052) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4371) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7222) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7466) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9959) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27395) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22430) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24236) * $signed(input_fmap_59[7:0]) +
	( 10'sd 269) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_61[7:0]) +
	( 13'sd 4055) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1195) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10218) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24360) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18205) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23080) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28861) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7540) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14586) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32735) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2996) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31523) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24468) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7688) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31892) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22470) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5971) * $signed(input_fmap_88[7:0]) +
	( 11'sd 656) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17371) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18029) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20683) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13797) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13389) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23295) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27434) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21454) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29329) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1253) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23467) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18251) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29180) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8927) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17603) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28619) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21368) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30912) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4957) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6575) * $signed(input_fmap_115[7:0]) +
	( 10'sd 321) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6395) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13862) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1472) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11761) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23757) * $signed(input_fmap_124[7:0]) +
	( 12'sd 2040) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17118) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_165;
assign conv_mac_165 = 
	( 16'sd 24232) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5762) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30629) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29421) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24133) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25093) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6457) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31075) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9466) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12157) * $signed(input_fmap_12[7:0]) +
	( 10'sd 378) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18492) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27897) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29685) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26381) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27044) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23289) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20743) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30964) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_24[7:0]) +
	( 9'sd 173) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1192) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13346) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7067) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12629) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25176) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25210) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19466) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3473) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6359) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26916) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6349) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1497) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8668) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23358) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10191) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23809) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26786) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20930) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28671) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12953) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21257) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18276) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24911) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18346) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12640) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32236) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24905) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27520) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7343) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22798) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26070) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25785) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2720) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_81[7:0]) +
	( 8'sd 65) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15316) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31800) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25807) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15036) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7572) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25976) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14089) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5576) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22834) * $signed(input_fmap_95[7:0]) +
	( 12'sd 2047) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26154) * $signed(input_fmap_98[7:0]) +
	( 5'sd 12) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12404) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13771) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6559) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24035) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3992) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30944) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10047) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9996) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24494) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17585) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27398) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17129) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14644) * $signed(input_fmap_117[7:0]) +
	( 10'sd 352) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15565) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26107) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24321) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3477) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_166;
assign conv_mac_166 = 
	( 15'sd 10467) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24158) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28433) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22501) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25859) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31219) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27543) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21469) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11218) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2501) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8130) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4641) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26392) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31259) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19584) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21909) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28648) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19605) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8771) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3830) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31464) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26895) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17039) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31595) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3642) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31603) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15070) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16337) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19089) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13506) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21212) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9122) * $signed(input_fmap_50[7:0]) +
	( 9'sd 205) * $signed(input_fmap_51[7:0]) +
	( 9'sd 206) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6969) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15778) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15425) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20006) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13120) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18332) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1220) * $signed(input_fmap_67[7:0]) +
	( 11'sd 976) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25949) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8846) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30419) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5364) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26449) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17990) * $signed(input_fmap_78[7:0]) +
	( 10'sd 386) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14892) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5711) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6265) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29776) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22397) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9491) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2809) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6319) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20402) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29320) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14000) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4459) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22282) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18976) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24235) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10989) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11292) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27774) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21126) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_108[7:0]) +
	( 14'sd 8118) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14614) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17359) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25677) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6069) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31005) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26207) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23365) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28038) * $signed(input_fmap_118[7:0]) +
	( 11'sd 579) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22191) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6709) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6516) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4626) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_167;
assign conv_mac_167 = 
	( 16'sd 18792) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11127) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30110) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8463) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_5[7:0]) +
	( 11'sd 741) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29680) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20683) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28395) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32762) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27123) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22900) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2479) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11666) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27872) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5729) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10414) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3042) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14522) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32484) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23094) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26730) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27760) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5879) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12087) * $signed(input_fmap_38[7:0]) +
	( 11'sd 623) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13308) * $signed(input_fmap_40[7:0]) +
	( 10'sd 393) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2557) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28296) * $signed(input_fmap_44[7:0]) +
	( 12'sd 2033) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20630) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1165) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24437) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20754) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11152) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17398) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14100) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30816) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23034) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5496) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16776) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21783) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31220) * $signed(input_fmap_67[7:0]) +
	( 9'sd 154) * $signed(input_fmap_68[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26867) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21100) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7477) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12210) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20162) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7841) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18233) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12736) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11488) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10423) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7195) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_91[7:0]) +
	( 11'sd 668) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2336) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27886) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9918) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5203) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10345) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18883) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26726) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6072) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25533) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19604) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27354) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6023) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_120[7:0]) +
	( 11'sd 735) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14275) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15042) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_168;
assign conv_mac_168 = 
	( 15'sd 13133) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16652) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19177) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18335) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9039) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30723) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17019) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25597) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25322) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3076) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6465) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20565) * $signed(input_fmap_23[7:0]) +
	( 11'sd 570) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21699) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18708) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13570) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13129) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27107) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32295) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20411) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26287) * $signed(input_fmap_34[7:0]) +
	( 11'sd 756) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27604) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6272) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27017) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30410) * $signed(input_fmap_40[7:0]) +
	( 9'sd 250) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6450) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7198) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5209) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17413) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16110) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10473) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25313) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9601) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10912) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1053) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16893) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25882) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20452) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18834) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9947) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20000) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30619) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31630) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15754) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7202) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9468) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1423) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17036) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9759) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18468) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20690) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18488) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28225) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13296) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_81[7:0]) +
	( 11'sd 881) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16600) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24427) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4674) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5448) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13528) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3973) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13433) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28704) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_100[7:0]) +
	( 11'sd 541) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24143) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17700) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28408) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14705) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32324) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9567) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31496) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6686) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22171) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7138) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12220) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8767) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22044) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_169;
assign conv_mac_169 = 
	( 16'sd 24394) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23841) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5144) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1951) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7842) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12658) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20644) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30290) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12943) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13615) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7837) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6895) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2961) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14932) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9719) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31935) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28648) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21327) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17896) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20156) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32689) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28430) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11119) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4628) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22602) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8197) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23722) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27689) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11104) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28494) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3613) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14510) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29983) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17223) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32247) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17735) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25438) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26910) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3432) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_54[7:0]) +
	( 11'sd 834) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26039) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22136) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13560) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16426) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20346) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3535) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10246) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7847) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32164) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7272) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8749) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16596) * $signed(input_fmap_76[7:0]) +
	( 12'sd 2027) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8973) * $signed(input_fmap_80[7:0]) +
	( 11'sd 1012) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18224) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30205) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16675) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18037) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11844) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21817) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27934) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28863) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16320) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18008) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3069) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12383) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18184) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_101[7:0]) +
	( 11'sd 714) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3246) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5182) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18882) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30231) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30144) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15272) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_110[7:0]) +
	( 7'sd 36) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27180) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8561) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31133) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18648) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23050) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7795) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16179) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30535) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18085) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21632) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16762) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_170;
assign conv_mac_170 = 
	( 14'sd 7035) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2595) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6528) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13061) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16636) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29060) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13979) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25870) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17920) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14034) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22914) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27104) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3809) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22722) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17018) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8709) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18301) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32489) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5056) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28493) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27401) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21619) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26705) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3873) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5538) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_40[7:0]) +
	( 13'sd 4024) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30551) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6455) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30286) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6657) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23503) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1960) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_51[7:0]) +
	( 10'sd 393) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25972) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23594) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31691) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29733) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30436) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22271) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3183) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3884) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21396) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29136) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16286) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15582) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12789) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31511) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6617) * $signed(input_fmap_72[7:0]) +
	( 11'sd 587) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23263) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22331) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21820) * $signed(input_fmap_76[7:0]) +
	( 10'sd 465) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24940) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19423) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17110) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5337) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8494) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18476) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28619) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8723) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30294) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25522) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16819) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13969) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21207) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24643) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26839) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26935) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1552) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13132) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23009) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15972) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16538) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27228) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20770) * $signed(input_fmap_115[7:0]) +
	( 11'sd 528) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5253) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31957) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21432) * $signed(input_fmap_126[7:0]) +
	( 12'sd 2045) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_171;
assign conv_mac_171 = 
	( 15'sd 10878) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18961) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29113) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30966) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11808) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8274) * $signed(input_fmap_11[7:0]) +
	( 11'sd 888) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21045) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20143) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17438) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12940) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27437) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17829) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3564) * $signed(input_fmap_23[7:0]) +
	( 11'sd 943) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11212) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18419) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17604) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17227) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18423) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5614) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2858) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17371) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1662) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28538) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13888) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16306) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15541) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14031) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21112) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20768) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10049) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_53[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7869) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17813) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25762) * $signed(input_fmap_57[7:0]) +
	( 11'sd 688) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11296) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21617) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_61[7:0]) +
	( 10'sd 358) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29003) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31935) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20522) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15015) * $signed(input_fmap_67[7:0]) +
	( 11'sd 899) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26168) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7243) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13790) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25413) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22659) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18336) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27873) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20340) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6451) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15993) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21029) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20092) * $signed(input_fmap_85[7:0]) +
	( 11'sd 745) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7084) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14351) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3640) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13073) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32410) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13469) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25735) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5258) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14412) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11854) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15445) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8320) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30604) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2095) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4144) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4161) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23474) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4503) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25636) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26938) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9713) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13812) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4606) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4589) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25986) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16210) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31534) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26248) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_172;
assign conv_mac_172 = 
	( 16'sd 18359) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31198) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22941) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9417) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11623) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26059) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9800) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25441) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18654) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1734) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22964) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24442) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12101) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_19[7:0]) +
	( 10'sd 375) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5697) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9136) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9478) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24892) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6663) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2498) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13598) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5764) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16073) * $signed(input_fmap_37[7:0]) +
	( 11'sd 730) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13411) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21692) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4375) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27072) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7986) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11481) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10081) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20737) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10620) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28149) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15153) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27458) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28212) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3550) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11925) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5964) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17680) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18985) * $signed(input_fmap_67[7:0]) +
	( 10'sd 352) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14194) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17863) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27918) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4105) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30518) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30360) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32643) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30297) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26495) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28192) * $signed(input_fmap_79[7:0]) +
	( 13'sd 4082) * $signed(input_fmap_80[7:0]) +
	( 6'sd 28) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21694) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17383) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17981) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26526) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8972) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8619) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12525) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4934) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29354) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8140) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21195) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29933) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11906) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16649) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19757) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8642) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25330) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28393) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14998) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14998) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19935) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31016) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29676) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27371) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16524) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11411) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4503) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1874) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_124[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4549) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_173;
assign conv_mac_173 = 
	( 15'sd 11141) * $signed(input_fmap_0[7:0]) +
	( 11'sd 1004) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23183) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24469) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13885) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7161) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15913) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28494) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31892) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9208) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21176) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17428) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30579) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21490) * $signed(input_fmap_23[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12293) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11223) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30618) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24931) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29086) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20253) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11622) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6619) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30506) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26311) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14154) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6231) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3638) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16357) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7241) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20509) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23587) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16468) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6285) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1828) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12400) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21984) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30522) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25579) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5742) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19454) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4468) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30594) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11576) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1687) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21215) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29334) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27435) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20858) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20392) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22607) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17175) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29999) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16774) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1625) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18005) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9121) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15304) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19724) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11588) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12958) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26748) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17324) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24844) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19604) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26061) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7598) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23763) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28898) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20150) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8223) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30932) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25937) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21791) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10807) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21100) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19080) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18122) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32256) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17247) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24506) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10421) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32262) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29500) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17315) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18492) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_174;
assign conv_mac_174 = 
	( 16'sd 29806) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28168) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32036) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6811) * $signed(input_fmap_5[7:0]) +
	( 10'sd 405) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16507) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30144) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14593) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18042) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10779) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10839) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_14[7:0]) +
	( 14'sd 8055) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28416) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15633) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18824) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_24[7:0]) +
	( 11'sd 653) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19560) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9663) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22851) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18832) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24560) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27841) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25708) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20142) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26783) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10864) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28114) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_43[7:0]) +
	( 11'sd 782) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22628) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21443) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17051) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25751) * $signed(input_fmap_48[7:0]) +
	( 8'sd 79) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24339) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22501) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15985) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6138) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3172) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20863) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25920) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12042) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3381) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_61[7:0]) +
	( 11'sd 781) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13226) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21921) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27276) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30651) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24831) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29384) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1390) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16690) * $signed(input_fmap_72[7:0]) +
	( 11'sd 873) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17494) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20788) * $signed(input_fmap_75[7:0]) +
	( 10'sd 492) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18557) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28199) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11358) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7808) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31043) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17691) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_96[7:0]) +
	( 10'sd 343) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31977) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13754) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13178) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27135) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27853) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7432) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10505) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9070) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26228) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28533) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12696) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9238) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19996) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9794) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13820) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11414) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23574) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10666) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18211) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1882) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32187) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22305) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_175;
assign conv_mac_175 = 
	( 14'sd 5385) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23801) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10132) * $signed(input_fmap_3[7:0]) +
	( 11'sd 899) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14153) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12726) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7505) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16767) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22171) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14751) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30087) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10357) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15040) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7283) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4781) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24159) * $signed(input_fmap_23[7:0]) +
	( 10'sd 379) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31261) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8450) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18881) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6824) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26625) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13550) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22283) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26406) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7629) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14164) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23161) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26955) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26300) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29973) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3426) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16495) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16483) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3143) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31524) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6111) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15288) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22947) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4226) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16425) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25040) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17149) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18214) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27674) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26570) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13217) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16913) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6466) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10207) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5302) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14926) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20050) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20668) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19011) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10865) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10257) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19926) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21829) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20766) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14401) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5827) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3827) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18949) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26983) * $signed(input_fmap_100[7:0]) +
	( 10'sd 494) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25216) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10788) * $signed(input_fmap_110[7:0]) +
	( 6'sd 25) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16659) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7864) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27521) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16230) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24703) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18884) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13075) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18988) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20667) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_176;
assign conv_mac_176 = 
	( 16'sd 25384) * $signed(input_fmap_0[7:0]) +
	( 7'sd 39) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14822) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5406) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30698) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26057) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2318) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13926) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26166) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17011) * $signed(input_fmap_16[7:0]) +
	( 12'sd 2026) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10316) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27456) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26390) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13475) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12959) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16545) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20934) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29245) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12927) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14854) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22711) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4676) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30429) * $signed(input_fmap_45[7:0]) +
	( 11'sd 1002) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6395) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31686) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14843) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13068) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17720) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31073) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31284) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17805) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26413) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11407) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18088) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26190) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_72[7:0]) +
	( 8'sd 104) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12821) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32236) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20562) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30933) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10811) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14490) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1734) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29287) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10947) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5195) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27822) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15635) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29662) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30608) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5829) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7774) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6384) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22931) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_102[7:0]) +
	( 11'sd 930) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19792) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28162) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11046) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16023) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15408) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5500) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25760) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4336) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11220) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31691) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28232) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4376) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15390) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31261) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16372) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_177;
assign conv_mac_177 = 
	( 16'sd 16582) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16747) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1399) * $signed(input_fmap_2[7:0]) +
	( 11'sd 630) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26102) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28838) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32687) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22078) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4658) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14567) * $signed(input_fmap_9[7:0]) +
	( 11'sd 752) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18246) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26904) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26962) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15238) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14293) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27147) * $signed(input_fmap_21[7:0]) +
	( 10'sd 493) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3934) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21675) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3671) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20793) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22039) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6983) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18282) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18362) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3679) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23345) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22007) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29424) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31278) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29853) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_42[7:0]) +
	( 11'sd 754) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13269) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27708) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8979) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18035) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5867) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18397) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11150) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4885) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21202) * $signed(input_fmap_55[7:0]) +
	( 11'sd 772) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27970) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18915) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32024) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24948) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23366) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29159) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27798) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19443) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17366) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19973) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26139) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21963) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25862) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18637) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19800) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15806) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16100) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23814) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13890) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12583) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20371) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7722) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4887) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16205) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8021) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19318) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29686) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8415) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9324) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27371) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32311) * $signed(input_fmap_101[7:0]) +
	( 11'sd 905) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18441) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11435) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22507) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26181) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16506) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5604) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26106) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21863) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2376) * $signed(input_fmap_116[7:0]) +
	( 10'sd 478) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16406) * $signed(input_fmap_118[7:0]) +
	( 10'sd 289) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16865) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_122[7:0]) +
	( 10'sd 272) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24895) * $signed(input_fmap_125[7:0]) +
	( 7'sd 61) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_178;
assign conv_mac_178 = 
	( 15'sd 13286) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7757) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23882) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9277) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1621) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26433) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28419) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12856) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17804) * $signed(input_fmap_19[7:0]) +
	( 11'sd 594) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2873) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19446) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13569) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26126) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21631) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29238) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19854) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14511) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18770) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17687) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19825) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2751) * $signed(input_fmap_37[7:0]) +
	( 11'sd 795) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24236) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10044) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23039) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16788) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24567) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12850) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3788) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30048) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13434) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5363) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10547) * $signed(input_fmap_55[7:0]) +
	( 11'sd 583) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1772) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10745) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30718) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9280) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20912) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10034) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15958) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20747) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15642) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26720) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4225) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1998) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21716) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15174) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7131) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19409) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23303) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21359) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12164) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1352) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30223) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19387) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15937) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3080) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6534) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14982) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15093) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11453) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3365) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15342) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8810) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17212) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23048) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29449) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16293) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32441) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12841) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17333) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4980) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29414) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26639) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21313) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10878) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11003) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_179;
assign conv_mac_179 = 
	( 15'sd 15219) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11291) * $signed(input_fmap_3[7:0]) +
	( 11'sd 607) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21088) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1966) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12936) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1407) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30349) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30245) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26502) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12623) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4479) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8114) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2729) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2085) * $signed(input_fmap_20[7:0]) +
	( 10'sd 301) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21161) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20714) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8775) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31330) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4774) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9191) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14753) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28476) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2982) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29155) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21040) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19873) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12549) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16212) * $signed(input_fmap_46[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31741) * $signed(input_fmap_48[7:0]) +
	( 14'sd 8163) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15189) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11958) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15866) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8959) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28124) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27192) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1324) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32070) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26102) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6765) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17039) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12211) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1877) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15133) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18720) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16310) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14764) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25850) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30149) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30064) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9614) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6919) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13035) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30059) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3973) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11080) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14028) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7009) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2467) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18202) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18835) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25924) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23068) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23886) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23628) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22308) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15381) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24339) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1142) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30215) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22822) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6550) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29507) * $signed(input_fmap_117[7:0]) +
	( 10'sd 387) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29996) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20541) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25715) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12221) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30225) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21688) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28707) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_180;
assign conv_mac_180 = 
	( 15'sd 14572) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10130) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27538) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10446) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24039) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9710) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24743) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1946) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15099) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28406) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19315) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10683) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4383) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28338) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30380) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13144) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18107) * $signed(input_fmap_21[7:0]) +
	( 10'sd 308) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19415) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10506) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31944) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31070) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28195) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27938) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21738) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22616) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9662) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25586) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31647) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14247) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28749) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7536) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18421) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20055) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2275) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9322) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11010) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26558) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29736) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10480) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24738) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12532) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18738) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25304) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11424) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20401) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7842) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5029) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3317) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25090) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9311) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32188) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25770) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12990) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3181) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4769) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26082) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30375) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29676) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18139) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24219) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2113) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5400) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25743) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23041) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23839) * $signed(input_fmap_95[7:0]) +
	( 7'sd 48) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22101) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16330) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26528) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28736) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21984) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23417) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24910) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17050) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27646) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7630) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17242) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27097) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12097) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26203) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17671) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32043) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22118) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19423) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28082) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30507) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_181;
assign conv_mac_181 = 
	( 16'sd 27993) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2105) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30319) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24754) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9925) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26055) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11595) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7858) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12040) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10055) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6992) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7757) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15873) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26078) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17696) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20649) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30064) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31973) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14114) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23308) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23147) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13294) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25017) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9778) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23262) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14727) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29708) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17646) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10733) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22789) * $signed(input_fmap_53[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8205) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12792) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17336) * $signed(input_fmap_59[7:0]) +
	( 10'sd 391) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28585) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30699) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8658) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24871) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4971) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_69[7:0]) +
	( 14'sd 8093) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20888) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27414) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_73[7:0]) +
	( 11'sd 1014) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20549) * $signed(input_fmap_76[7:0]) +
	( 11'sd 980) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8489) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11260) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31435) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27356) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11180) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3644) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28399) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14856) * $signed(input_fmap_96[7:0]) +
	( 10'sd 389) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2247) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28585) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16393) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9294) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10526) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31777) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15357) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27184) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29206) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22305) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16937) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22931) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24026) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4174) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3132) * $signed(input_fmap_125[7:0]) +
	( 11'sd 698) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3385) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_182;
assign conv_mac_182 = 
	( 16'sd 26765) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8410) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8760) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5350) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31864) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23838) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22495) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28368) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16616) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17595) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3800) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9752) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26183) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17149) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8974) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17115) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3881) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15358) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_32[7:0]) +
	( 8'sd 86) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6401) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11706) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22508) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25742) * $signed(input_fmap_38[7:0]) +
	( 11'sd 975) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4715) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11039) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15382) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26963) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22581) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25609) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25082) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4427) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29259) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24305) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15599) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11436) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19463) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22977) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14208) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25035) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4725) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11728) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4718) * $signed(input_fmap_67[7:0]) +
	( 14'sd 8163) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28379) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10391) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21655) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27409) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8382) * $signed(input_fmap_76[7:0]) +
	( 11'sd 907) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12980) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29825) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29609) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1185) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_82[7:0]) +
	( 11'sd 958) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30222) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16429) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23952) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8759) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5682) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11812) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7861) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25107) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1976) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23830) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14598) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22363) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10995) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4248) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29308) * $signed(input_fmap_118[7:0]) +
	( 13'sd 4008) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4306) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22424) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17248) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12969) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7355) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_183;
assign conv_mac_183 = 
	( 16'sd 17416) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5999) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24432) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30225) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3924) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29717) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19764) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15689) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26025) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22435) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20550) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17786) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27314) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21149) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25634) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21062) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27343) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16333) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15986) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5324) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13578) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24945) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30502) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16962) * $signed(input_fmap_40[7:0]) +
	( 11'sd 655) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6180) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10249) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4725) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2451) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_46[7:0]) +
	( 11'sd 971) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3313) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10471) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7839) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12722) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28870) * $signed(input_fmap_58[7:0]) +
	( 7'sd 51) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29253) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1964) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32045) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4411) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31475) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1434) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29487) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7858) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11110) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1215) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30191) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_78[7:0]) +
	( 10'sd 428) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17971) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27857) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16194) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31327) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29216) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3626) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3265) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26508) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6595) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22101) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12107) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19126) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6509) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26094) * $signed(input_fmap_97[7:0]) +
	( 8'sd 82) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17953) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14336) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13704) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4928) * $signed(input_fmap_102[7:0]) +
	( 11'sd 792) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21530) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1706) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5088) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23036) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16976) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24506) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28579) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29634) * $signed(input_fmap_117[7:0]) +
	( 11'sd 682) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8970) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24702) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26806) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31989) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30568) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30552) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_184;
assign conv_mac_184 = 
	( 15'sd 15628) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18981) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20316) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19615) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3458) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14742) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9220) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2873) * $signed(input_fmap_13[7:0]) +
	( 10'sd 415) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21335) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31427) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7524) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2094) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7251) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5784) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3659) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27609) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_31[7:0]) +
	( 11'sd 632) * $signed(input_fmap_32[7:0]) +
	( 11'sd 632) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_37[7:0]) +
	( 7'sd 32) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20359) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24188) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22679) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14516) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30577) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5236) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13019) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20307) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19965) * $signed(input_fmap_50[7:0]) +
	( 15'sd 16215) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6160) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20506) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30105) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13479) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25435) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24140) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23731) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4406) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6721) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21429) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20167) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21736) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13375) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14236) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32077) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26541) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26714) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7756) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9678) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11373) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25495) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26738) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2495) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31329) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29283) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9732) * $signed(input_fmap_88[7:0]) +
	( 9'sd 129) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31388) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23863) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10136) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21279) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25227) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25647) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2152) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20065) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20035) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3264) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17819) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13354) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2248) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7070) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8436) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31588) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17955) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18591) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9569) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15271) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25489) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31426) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4252) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13874) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_123[7:0]) +
	( 11'sd 991) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5618) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16687) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_185;
assign conv_mac_185 = 
	( 10'sd 263) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25846) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10609) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6860) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18344) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21993) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_10[7:0]) +
	( 7'sd 36) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7125) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5468) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30373) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28765) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18840) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20330) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26116) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2567) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21185) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17793) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11436) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18989) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30051) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22143) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17272) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8627) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4747) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17580) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27400) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6308) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12277) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9498) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20490) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32491) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20593) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19275) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29439) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15561) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20784) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27987) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7495) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25199) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27225) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27618) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28969) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31730) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11029) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21433) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23450) * $signed(input_fmap_86[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24607) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17675) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14460) * $signed(input_fmap_91[7:0]) +
	( 11'sd 842) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3164) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22870) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21845) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27871) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22697) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22636) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28279) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31243) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15642) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18533) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26644) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2771) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24960) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5050) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26130) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5695) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26037) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2959) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19893) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21509) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5439) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21561) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17845) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_186;
assign conv_mac_186 = 
	( 13'sd 2871) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22503) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31117) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13177) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_10[7:0]) +
	( 9'sd 192) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3485) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13348) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19257) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1869) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8318) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1867) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9511) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30967) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25605) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15828) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31551) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24144) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6519) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3988) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12493) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5417) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19966) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11296) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32743) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28876) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8273) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31509) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16987) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12317) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3806) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22207) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18487) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26373) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7995) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20779) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22505) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14284) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17439) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28745) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18298) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3469) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26189) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6107) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22263) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6794) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24981) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23172) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16027) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31528) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26204) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11915) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17248) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24610) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1874) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6519) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32488) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23384) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30272) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21166) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4545) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25618) * $signed(input_fmap_99[7:0]) +
	( 10'sd 354) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13524) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11173) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2147) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_107[7:0]) +
	( 5'sd 13) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27154) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21264) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27273) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5547) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11535) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25430) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31943) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26542) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30346) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23035) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_187;
assign conv_mac_187 = 
	( 15'sd 10501) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17400) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9174) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11008) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4732) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15370) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6728) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6163) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21375) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7106) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8893) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18549) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17969) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10885) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17916) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18282) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12148) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17023) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32442) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_27[7:0]) +
	( 9'sd 130) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29632) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5328) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6906) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9686) * $signed(input_fmap_32[7:0]) +
	( 10'sd 426) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23290) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28865) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14988) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17618) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19787) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29605) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30410) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11886) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_48[7:0]) +
	( 11'sd 972) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9608) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7643) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10238) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10665) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20188) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31815) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18758) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5677) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9719) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24524) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4213) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11302) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30873) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20127) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20246) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11119) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8743) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13169) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26746) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24481) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9801) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31669) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19816) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2921) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18970) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22389) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21176) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_84[7:0]) +
	( 11'sd 813) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15418) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2639) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15370) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13561) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11884) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16747) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21796) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30147) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1997) * $signed(input_fmap_97[7:0]) +
	( 11'sd 713) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1109) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3251) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23365) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11568) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4456) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20658) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9686) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26312) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3855) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12833) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23087) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19362) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18207) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14422) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18060) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24688) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14189) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_188;
assign conv_mac_188 = 
	( 16'sd 26617) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28159) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3174) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5798) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18253) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20220) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26145) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2580) * $signed(input_fmap_9[7:0]) +
	( 10'sd 282) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11439) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10374) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17602) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32558) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7584) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32504) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6756) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30137) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29024) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27511) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15669) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14921) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28775) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5379) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29721) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19925) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1505) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20000) * $signed(input_fmap_37[7:0]) +
	( 10'sd 419) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6695) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6000) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29446) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30157) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24659) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23637) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9356) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15515) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15340) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30209) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5151) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17102) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1781) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23412) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22000) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30882) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16038) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24617) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23159) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8281) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12206) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19583) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22807) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4629) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31363) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1306) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11111) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2915) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27418) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1994) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25573) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7703) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11065) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9003) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7160) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5689) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5020) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13041) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9488) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31152) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28967) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17895) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22264) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9137) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7342) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22936) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28115) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30086) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18123) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11263) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6556) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21640) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31336) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24108) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6839) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21532) * $signed(input_fmap_119[7:0]) +
	( 11'sd 517) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2727) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18888) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23843) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_189;
assign conv_mac_189 = 
	( 12'sd 1037) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11865) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19236) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25143) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24533) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12016) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29434) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12995) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10989) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13306) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7803) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14889) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9622) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22562) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1729) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29753) * $signed(input_fmap_32[7:0]) +
	( 10'sd 393) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10794) * $signed(input_fmap_34[7:0]) +
	( 11'sd 935) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3214) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31219) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22375) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3835) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15617) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7771) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1488) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14294) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13481) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20720) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24174) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3925) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24362) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3728) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21305) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24867) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22977) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6420) * $signed(input_fmap_66[7:0]) +
	( 10'sd 472) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16935) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31011) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4151) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6383) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18594) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18532) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12719) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6377) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15608) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21459) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14326) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9282) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21005) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18132) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1440) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26148) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31602) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20936) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25129) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28767) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8442) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1486) * $signed(input_fmap_106[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2990) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20953) * $signed(input_fmap_111[7:0]) +
	( 13'sd 4075) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25276) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14441) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21060) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18955) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8634) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4486) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26003) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28694) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_190;
assign conv_mac_190 = 
	( 14'sd 5378) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9185) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22552) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20977) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11991) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3417) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16263) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28960) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9966) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30998) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12733) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29433) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1284) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21034) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25761) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18945) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15573) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26685) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4205) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5717) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9348) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2434) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28976) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26465) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4935) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8608) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29632) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_39[7:0]) +
	( 11'sd 983) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2379) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12358) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19029) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27018) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7309) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14746) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28268) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2680) * $signed(input_fmap_52[7:0]) +
	( 9'sd 193) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1623) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27634) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11200) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25799) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4576) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10075) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16780) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20440) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30881) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8379) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9192) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24063) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30108) * $signed(input_fmap_74[7:0]) +
	( 11'sd 529) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14625) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2790) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29869) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8620) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20494) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5085) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28173) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6014) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1677) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20561) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_97[7:0]) +
	( 10'sd 257) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17927) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4346) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8223) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29311) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13144) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21454) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13680) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7606) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25500) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7618) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19030) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20846) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18721) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15559) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14412) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2745) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27422) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31675) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23340) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_191;
assign conv_mac_191 = 
	( 16'sd 16461) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1518) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9840) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30050) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16147) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18203) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14056) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31922) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24560) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6932) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19784) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29055) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25755) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28453) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17115) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23666) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26190) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1566) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17543) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31831) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26382) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19966) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6672) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20518) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12548) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5220) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19658) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23538) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29605) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3846) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13621) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1181) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32482) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8534) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25328) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3456) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14984) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31448) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31498) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20620) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9899) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25901) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28761) * $signed(input_fmap_56[7:0]) +
	( 11'sd 758) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20615) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8283) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32754) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11961) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30529) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31200) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28267) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17752) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5751) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18649) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32721) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11758) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9855) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31974) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7475) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24316) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29949) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22304) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27274) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22705) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29101) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32667) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25419) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32512) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25805) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5708) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8535) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29945) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13423) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23805) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9142) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21968) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25072) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3417) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29428) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26995) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25035) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16661) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9543) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_192;
assign conv_mac_192 = 
	( 16'sd 25516) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19502) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32764) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23011) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6333) * $signed(input_fmap_4[7:0]) +
	( 11'sd 697) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15177) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29549) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18704) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14082) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17973) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19883) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12117) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4583) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12177) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7423) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5678) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6776) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15203) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27103) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8471) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10453) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29116) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9321) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4649) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26901) * $signed(input_fmap_40[7:0]) +
	( 11'sd 839) * $signed(input_fmap_41[7:0]) +
	( 11'sd 523) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_43[7:0]) +
	( 11'sd 835) * $signed(input_fmap_44[7:0]) +
	( 11'sd 974) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22302) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_47[7:0]) +
	( 7'sd 41) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6881) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11094) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12797) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5029) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22534) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2785) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7085) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_58[7:0]) +
	( 9'sd 194) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2052) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6040) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29320) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1709) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4611) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21826) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9740) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25189) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20933) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16275) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30500) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18504) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2471) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30368) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10076) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2859) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15203) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8944) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23755) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6616) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25300) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29313) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14586) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16346) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31361) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17918) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17819) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6341) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22952) * $signed(input_fmap_101[7:0]) +
	( 9'sd 180) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21869) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27095) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32285) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31537) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20877) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11133) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10364) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18604) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32226) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2846) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1134) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31947) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27095) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26605) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30494) * $signed(input_fmap_126[7:0]) +
	( 11'sd 979) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_193;
assign conv_mac_193 = 
	( 16'sd 22405) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6122) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23938) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15483) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3514) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21651) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6596) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2564) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15555) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22317) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8900) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20142) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30956) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23581) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10081) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5315) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9460) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22875) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9408) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14928) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10501) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23693) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14967) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28714) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23924) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15564) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22065) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22023) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21480) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4545) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13676) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30447) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8210) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11573) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29377) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18307) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26209) * $signed(input_fmap_59[7:0]) +
	( 11'sd 974) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11407) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27540) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26977) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19962) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18284) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13290) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15975) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8202) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17474) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25986) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27736) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15330) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2317) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1712) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27965) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31037) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21185) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4100) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8982) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19354) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16381) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26968) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12233) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23612) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30544) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26886) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7049) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24276) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2681) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12345) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13668) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2471) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11580) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22702) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1233) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28644) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26054) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4301) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26946) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16818) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9324) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24286) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_194;
assign conv_mac_194 = 
	( 16'sd 21126) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27150) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31058) * $signed(input_fmap_4[7:0]) +
	( 10'sd 336) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3334) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26966) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25264) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8386) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7897) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18918) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22455) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28261) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5172) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23738) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10535) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28947) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21189) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16781) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2433) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15568) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13409) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13714) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4629) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27137) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1353) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9554) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29170) * $signed(input_fmap_45[7:0]) +
	( 11'sd 839) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2280) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13113) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23576) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28937) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13314) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14671) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30629) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16428) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24960) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18283) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20308) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2500) * $signed(input_fmap_64[7:0]) +
	( 11'sd 619) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19428) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15537) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_68[7:0]) +
	( 11'sd 936) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26285) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3796) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15415) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8979) * $signed(input_fmap_74[7:0]) +
	( 14'sd 8139) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17721) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10912) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7313) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10884) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5006) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16497) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20606) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12951) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14364) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5086) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32499) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29638) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25799) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1264) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13795) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25314) * $signed(input_fmap_100[7:0]) +
	( 10'sd 325) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12050) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21489) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28177) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24442) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5253) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29776) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6997) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8407) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11145) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12880) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25507) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25585) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28742) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29630) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15846) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10283) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2597) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_195;
assign conv_mac_195 = 
	( 16'sd 22392) * $signed(input_fmap_0[7:0]) +
	( 11'sd 848) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3143) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1789) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2071) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10817) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3776) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29746) * $signed(input_fmap_16[7:0]) +
	( 11'sd 682) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24549) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18301) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_20[7:0]) +
	( 10'sd 294) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7719) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18387) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10502) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17387) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16775) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5960) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21303) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22614) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7162) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11585) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4886) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29951) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26758) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16826) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21720) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19206) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8775) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17546) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7318) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28537) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3780) * $signed(input_fmap_51[7:0]) +
	( 11'sd 602) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27733) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28753) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23669) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9788) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27353) * $signed(input_fmap_65[7:0]) +
	( 11'sd 542) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13318) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20738) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5550) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14689) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13105) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18749) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21080) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11230) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28843) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20870) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12540) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24100) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3266) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29053) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17215) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24007) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26029) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29556) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14717) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26652) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14349) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6794) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18095) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6051) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26637) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17746) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24728) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32062) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18053) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7942) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5914) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32035) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22414) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24760) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17429) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20166) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22848) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19358) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8255) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11477) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20745) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_196;
assign conv_mac_196 = 
	( 16'sd 16682) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28636) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_3[7:0]) +
	( 9'sd 232) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32365) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30959) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11461) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24322) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17964) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5875) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22910) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7711) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26441) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11237) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30118) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10762) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31904) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5957) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31209) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15701) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27466) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12586) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8734) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21641) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16429) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12995) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15261) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32432) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7351) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22768) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1459) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31061) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19128) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8913) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26076) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27453) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9097) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16310) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13745) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9370) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7711) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4103) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18097) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21357) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27961) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25532) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2325) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12263) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17869) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17809) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25885) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5151) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30958) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3448) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5697) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28321) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26741) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7494) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13043) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1154) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29436) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7793) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26160) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3453) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3990) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15082) * $signed(input_fmap_90[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2270) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5787) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27902) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25631) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22519) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10911) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14381) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31191) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9533) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12655) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27605) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30689) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28368) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15566) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9486) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9030) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15235) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10373) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14072) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29936) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_197;
assign conv_mac_197 = 
	( 15'sd 11039) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_1[7:0]) +
	( 11'sd 609) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15262) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4935) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29969) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14617) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9586) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5590) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22176) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19330) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32167) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29837) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30968) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19404) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3275) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12536) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11283) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16061) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16167) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27160) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3880) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28484) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6109) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9654) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9751) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24569) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1459) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25295) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16800) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24127) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7588) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3045) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13629) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2392) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19383) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30628) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16887) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18807) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28546) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27730) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3920) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32004) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16167) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4158) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20901) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24662) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17731) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32214) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21037) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13003) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29912) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32214) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10469) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6059) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22270) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28770) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27383) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16145) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27628) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13211) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10017) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29571) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18258) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21185) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28634) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8153) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27440) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21756) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19409) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29215) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32403) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23114) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23178) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20436) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30753) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21406) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11150) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25433) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14253) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24950) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28506) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16207) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25399) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32034) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19822) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12257) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10976) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22504) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11576) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6457) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31671) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27739) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_198;
assign conv_mac_198 = 
	( 15'sd 13618) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15094) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6924) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11312) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32642) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19073) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2848) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12691) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18039) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5292) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28075) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5784) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26616) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12819) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16750) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21894) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12951) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12154) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14938) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31105) * $signed(input_fmap_25[7:0]) +
	( 10'sd 415) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3911) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32528) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11844) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19926) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23940) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6014) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10743) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14329) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25360) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24804) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11495) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26250) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12658) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18495) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15718) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12596) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4183) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25931) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8950) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17760) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21141) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20376) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22509) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28501) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28045) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5325) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19674) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21395) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16170) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19364) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14614) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12968) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22364) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9289) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10047) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8601) * $signed(input_fmap_81[7:0]) +
	( 10'sd 356) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26604) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2257) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16922) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5288) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14599) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25201) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24894) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12783) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24835) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19156) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3457) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9307) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31253) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7094) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10889) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13981) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22956) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11972) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23434) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28522) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24183) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21982) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31713) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28264) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6785) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15826) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10682) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_199;
assign conv_mac_199 = 
	( 15'sd 8721) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12165) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4353) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22260) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14113) * $signed(input_fmap_6[7:0]) +
	( 9'sd 220) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30315) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26285) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7512) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9634) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11940) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26450) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29259) * $signed(input_fmap_19[7:0]) +
	( 14'sd 8139) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26069) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30488) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4155) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19388) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6658) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23421) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13116) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25883) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14019) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23818) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11599) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7073) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12142) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4515) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3132) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12323) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9702) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6371) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16622) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6215) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26516) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28625) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30762) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6268) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20565) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7310) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7515) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2989) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16117) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16697) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32533) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27728) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26972) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3334) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31442) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7716) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29841) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4709) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30890) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19826) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15210) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22779) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12040) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31833) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4576) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3077) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6618) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32289) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17801) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18109) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11897) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28519) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7845) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20503) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3230) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31628) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5251) * $signed(input_fmap_112[7:0]) +
	( 11'sd 945) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25971) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2603) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10426) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5351) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3903) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8773) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12864) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18325) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_200;
assign conv_mac_200 = 
	( 16'sd 20767) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13286) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15823) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27609) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9481) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16771) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1381) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16198) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6258) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22457) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10449) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11445) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20007) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24995) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18029) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27483) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23816) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19129) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28084) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27339) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5036) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19145) * $signed(input_fmap_36[7:0]) +
	( 10'sd 428) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18880) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8876) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15617) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11166) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24503) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_45[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6257) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30311) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9801) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25339) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27882) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28633) * $signed(input_fmap_54[7:0]) +
	( 8'sd 89) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27108) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9359) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7986) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16596) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6520) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3579) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4930) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30689) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_71[7:0]) +
	( 11'sd 761) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13219) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24767) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11664) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17606) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1380) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9953) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4655) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20042) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1062) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23895) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10786) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15830) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15863) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22130) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4532) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16764) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11690) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28137) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15598) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29778) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8824) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30856) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14227) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1325) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3659) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5239) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20677) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11928) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22697) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26910) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27891) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22038) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8148) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21078) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18959) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29693) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16610) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_201;
assign conv_mac_201 = 
	( 16'sd 31980) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12260) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31127) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25905) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14189) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12139) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12448) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14500) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28182) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29530) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30974) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30583) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23170) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21532) * $signed(input_fmap_18[7:0]) +
	( 11'sd 869) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15018) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31144) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32448) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10635) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23689) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1121) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10799) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10417) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13676) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_36[7:0]) +
	( 11'sd 718) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_40[7:0]) +
	( 10'sd 325) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23990) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16261) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1618) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28641) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9415) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1341) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8028) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_55[7:0]) +
	( 11'sd 889) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15719) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32697) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7755) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30349) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14200) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30900) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32113) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32119) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17429) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25636) * $signed(input_fmap_71[7:0]) +
	( 11'sd 911) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21096) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29354) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24807) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22224) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28334) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9267) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17785) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13673) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28776) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10046) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5174) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20008) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23747) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9082) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21904) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22729) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20347) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22579) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23746) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20758) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_117[7:0]) +
	( 11'sd 642) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13488) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32488) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19356) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8890) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22831) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2341) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_202;
assign conv_mac_202 = 
	( 15'sd 15193) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12858) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7386) * $signed(input_fmap_3[7:0]) +
	( 11'sd 518) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27540) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19751) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23253) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16309) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2267) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5192) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7663) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5595) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19875) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31957) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9037) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3064) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2443) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14289) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32174) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18956) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13750) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25952) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20677) * $signed(input_fmap_40[7:0]) +
	( 14'sd 8055) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20906) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_43[7:0]) +
	( 9'sd 197) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31649) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20264) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16394) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21288) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29792) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27512) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15533) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9871) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28120) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31769) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22248) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3753) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1780) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26161) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9657) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21439) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10573) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23829) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9802) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30997) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18010) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30743) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13394) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22346) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14393) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13035) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2763) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6270) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16369) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2291) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7199) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5363) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19590) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1209) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17993) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18490) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18449) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_95[7:0]) +
	( 7'sd 53) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6574) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20948) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29392) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16832) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1059) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25045) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20963) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11187) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18575) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28288) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3438) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11808) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31711) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8981) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4100) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28294) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31699) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24396) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26477) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21754) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24732) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5933) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_203;
assign conv_mac_203 = 
	( 16'sd 19236) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28472) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12674) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20141) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26954) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4920) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1913) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28548) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2386) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_15[7:0]) +
	( 10'sd 379) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12530) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7398) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20851) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31853) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_24[7:0]) +
	( 11'sd 548) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16692) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8623) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31237) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24157) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17061) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21423) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26448) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29293) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3179) * $signed(input_fmap_40[7:0]) +
	( 11'sd 997) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4617) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13307) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_45[7:0]) +
	( 11'sd 721) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26307) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19958) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18370) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12635) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6694) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9031) * $signed(input_fmap_53[7:0]) +
	( 11'sd 571) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4503) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15130) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24013) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16681) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8365) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23639) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30599) * $signed(input_fmap_63[7:0]) +
	( 11'sd 536) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28298) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10682) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14712) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30793) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21547) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7295) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25877) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_78[7:0]) +
	( 12'sd 2025) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7993) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_81[7:0]) +
	( 9'sd 134) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13187) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20216) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2082) * $signed(input_fmap_85[7:0]) +
	( 10'sd 262) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24629) * $signed(input_fmap_87[7:0]) +
	( 10'sd 274) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5965) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_90[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17216) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25667) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9204) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9547) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14299) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32072) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2226) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5645) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29032) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23704) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12450) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24874) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28694) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12416) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17336) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18356) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10303) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21926) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27425) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6705) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17777) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12715) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15974) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13626) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_204;
assign conv_mac_204 = 
	( 13'sd 3623) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31158) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25304) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2741) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10167) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16627) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17632) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16846) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24284) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1961) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21293) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14563) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26238) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11261) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31156) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4867) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4387) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20913) * $signed(input_fmap_25[7:0]) +
	( 11'sd 929) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4627) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10875) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22265) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7272) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24295) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23608) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26001) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22581) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27872) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26976) * $signed(input_fmap_39[7:0]) +
	( 11'sd 651) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30239) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19007) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31920) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1481) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6208) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3367) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12006) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12498) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9807) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25752) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15025) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18174) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19151) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15465) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5990) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17547) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8881) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32138) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28705) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_75[7:0]) +
	( 11'sd 592) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7276) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18733) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20899) * $signed(input_fmap_83[7:0]) +
	( 9'sd 160) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3802) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13530) * $signed(input_fmap_86[7:0]) +
	( 11'sd 953) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30346) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5761) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22360) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25268) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21068) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20642) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20938) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3011) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15975) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18678) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32450) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15573) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30953) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13165) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30423) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17914) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12795) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7970) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24259) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9855) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7458) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1590) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12435) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13184) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_205;
assign conv_mac_205 = 
	( 16'sd 28130) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18098) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10775) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22364) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27913) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25429) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27921) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31093) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17870) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3446) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28777) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24432) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6862) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31965) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20177) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25028) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32159) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27797) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18981) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2488) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19406) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20613) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9827) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2719) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18913) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1546) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31165) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9280) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6670) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19205) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26694) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4624) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19585) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20768) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31107) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30499) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21969) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6446) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4780) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27773) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1941) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23305) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32235) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_88[7:0]) +
	( 11'sd 774) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27685) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18854) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8233) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21456) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19225) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14352) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30055) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9038) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3003) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32232) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6908) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24725) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21969) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8868) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20167) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13711) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16155) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28185) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6694) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19604) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25400) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15650) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28799) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4363) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7140) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20828) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_206;
assign conv_mac_206 = 
	( 16'sd 23593) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17389) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19617) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7704) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1383) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30262) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_10[7:0]) +
	( 11'sd 535) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5943) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24942) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32145) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25424) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2543) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23623) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24722) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21430) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24615) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1950) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31896) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3521) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21336) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23110) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11122) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26150) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5883) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12305) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16596) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16887) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5700) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9486) * $signed(input_fmap_50[7:0]) +
	( 11'sd 687) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26119) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17493) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31636) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25224) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5199) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21245) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15798) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11915) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4831) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23364) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3660) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5267) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19344) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19234) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3770) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8506) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17911) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5623) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10327) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23034) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16407) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15732) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_85[7:0]) +
	( 10'sd 341) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3045) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2250) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8465) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17102) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22242) * $signed(input_fmap_93[7:0]) +
	( 11'sd 736) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19230) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6356) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18999) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28550) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21326) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20256) * $signed(input_fmap_103[7:0]) +
	( 10'sd 355) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12310) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13006) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4526) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32359) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7437) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7625) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18394) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3014) * $signed(input_fmap_115[7:0]) +
	( 11'sd 803) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1537) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25452) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28947) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27558) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15137) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18421) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_207;
assign conv_mac_207 = 
	( 14'sd 7353) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30326) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19243) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9831) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30500) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29192) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17779) * $signed(input_fmap_10[7:0]) +
	( 11'sd 714) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11882) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19275) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31032) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12956) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14597) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12023) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29317) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8274) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2160) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17355) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_27[7:0]) +
	( 10'sd 451) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6578) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16612) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1754) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19233) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20004) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2359) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21102) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1215) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28984) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24925) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29789) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11570) * $signed(input_fmap_44[7:0]) +
	( 11'sd 1013) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22704) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21479) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9435) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27023) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20057) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16180) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29383) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10683) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29397) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27909) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26727) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19641) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26349) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10215) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_71[7:0]) +
	( 10'sd 423) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23337) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31940) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24980) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27257) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24936) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11621) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30745) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1360) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21085) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2141) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26451) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7834) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_89[7:0]) +
	( 11'sd 729) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27514) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28731) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17046) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8705) * $signed(input_fmap_98[7:0]) +
	( 9'sd 221) * $signed(input_fmap_99[7:0]) +
	( 13'sd 4050) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22915) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13842) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18294) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28524) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_107[7:0]) +
	( 13'sd 4032) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10131) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18884) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16566) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31132) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24545) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4517) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23802) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21495) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18547) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24433) * $signed(input_fmap_118[7:0]) +
	( 11'sd 660) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29679) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26639) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9564) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28543) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20355) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20374) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_208;
assign conv_mac_208 = 
	( 15'sd 15640) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29944) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12659) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9748) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13344) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19015) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16043) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24831) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29303) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21167) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17104) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24442) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15293) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6698) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24874) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23209) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_28[7:0]) +
	( 10'sd 416) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32080) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19777) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32553) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32365) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28209) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25793) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30332) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17783) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19648) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1684) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30418) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_49[7:0]) +
	( 12'sd 2025) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20557) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18678) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12442) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20873) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5878) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18570) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9079) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13416) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29571) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22311) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16228) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3441) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10039) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25616) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26194) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28568) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19417) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30364) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8335) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16396) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28304) * $signed(input_fmap_83[7:0]) +
	( 10'sd 296) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19979) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19079) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27862) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3151) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5407) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31507) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14091) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30141) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23616) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9190) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12693) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16215) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22169) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24095) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26384) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16363) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22334) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21496) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17167) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5481) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7221) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15329) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15959) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19055) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7697) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_209;
assign conv_mac_209 = 
	( 15'sd 13712) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9119) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8611) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4179) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3424) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1192) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19802) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24811) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27146) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13544) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7169) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9771) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27321) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_25[7:0]) +
	( 10'sd 409) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25982) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22027) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7593) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5138) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30576) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5400) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30957) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12245) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3137) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28972) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27907) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8316) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32148) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31034) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31905) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25099) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6130) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17428) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21716) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31466) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12639) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30200) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21994) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22807) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4906) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9216) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22295) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14792) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6854) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22035) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14818) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4391) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5715) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21303) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11960) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24788) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28393) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17058) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9693) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22833) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32627) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12617) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2509) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4233) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22154) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27115) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26709) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30756) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19186) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29703) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9756) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30876) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25296) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12277) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29437) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22331) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15501) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14848) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25479) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17007) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11167) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19376) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22773) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_210;
assign conv_mac_210 = 
	( 16'sd 24966) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18635) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19172) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12985) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3664) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3320) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25513) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31538) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18826) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23377) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22888) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4942) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31001) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26135) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2456) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26430) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23578) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26928) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19168) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15046) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12941) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6802) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21192) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26350) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9765) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22324) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18934) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29028) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23013) * $signed(input_fmap_41[7:0]) +
	( 10'sd 268) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14656) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20313) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21135) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7905) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5380) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22575) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8643) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9673) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11649) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8981) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_55[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7065) * $signed(input_fmap_57[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32419) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9006) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10425) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_64[7:0]) +
	( 11'sd 941) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8240) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31764) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14526) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14355) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2236) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26624) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16776) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32682) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29576) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29921) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17304) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30119) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20279) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21276) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18328) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12320) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32732) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7536) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18467) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5319) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9830) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32726) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25957) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9052) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22007) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23429) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19361) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3232) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15978) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31955) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32121) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24385) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10210) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7355) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14528) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20502) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8469) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28141) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12402) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_211;
assign conv_mac_211 = 
	( 16'sd 24715) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30752) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22450) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11578) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14108) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10424) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10092) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29259) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23469) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16080) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10823) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26638) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10926) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7376) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7324) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19544) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18701) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16397) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15957) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21242) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27916) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13183) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3333) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12556) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32564) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19363) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6122) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2832) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4102) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4775) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31709) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22332) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6231) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12138) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24135) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20726) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_57[7:0]) +
	( 10'sd 458) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24272) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10131) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22960) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31047) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21648) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7048) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16268) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15729) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22727) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11061) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6673) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27876) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13614) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17762) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_77[7:0]) +
	( 11'sd 893) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_79[7:0]) +
	( 5'sd 8) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10882) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9849) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23121) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12648) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1657) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21726) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25623) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7398) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3695) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7827) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17109) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25818) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29623) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14526) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10407) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16189) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10097) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4807) * $signed(input_fmap_106[7:0]) +
	( 10'sd 285) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31116) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19842) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5413) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5851) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25084) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14435) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14152) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6317) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12286) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18496) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31650) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10024) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9561) * $signed(input_fmap_124[7:0]) +
	( 12'sd 2011) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1547) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1060) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_212;
assign conv_mac_212 = 
	( 16'sd 25347) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26479) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1466) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12492) * $signed(input_fmap_5[7:0]) +
	( 11'sd 516) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30774) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_9[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27390) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25736) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15115) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13889) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8578) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4187) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19177) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16873) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18424) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7558) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14155) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31043) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14836) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26109) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10255) * $signed(input_fmap_34[7:0]) +
	( 11'sd 873) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8833) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30029) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5656) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23503) * $signed(input_fmap_41[7:0]) +
	( 8'sd 70) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31624) * $signed(input_fmap_44[7:0]) +
	( 10'sd 316) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10470) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30944) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13452) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9697) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25320) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18809) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30701) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5665) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11205) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20519) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19388) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12292) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17046) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7147) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20049) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12902) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6249) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30121) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6504) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17876) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23577) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23855) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13228) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15980) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17944) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17052) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20015) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2339) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19940) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2817) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5136) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7524) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3742) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26926) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15797) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9985) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3177) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21440) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15331) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30885) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26682) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28960) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18871) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8319) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22445) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25515) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5686) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4893) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1974) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22127) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1518) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12274) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14776) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29253) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_213;
assign conv_mac_213 = 
	( 16'sd 25568) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18052) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32292) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26777) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31425) * $signed(input_fmap_7[7:0]) +
	( 13'sd 4028) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23343) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20456) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28083) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20895) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23394) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19425) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19366) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24786) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20403) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31358) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7873) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8106) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13677) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2096) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14427) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31577) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10169) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9581) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3547) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23119) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13487) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_43[7:0]) +
	( 7'sd 34) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2500) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26641) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25198) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8886) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11386) * $signed(input_fmap_52[7:0]) +
	( 11'sd 787) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_54[7:0]) +
	( 11'sd 773) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10333) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10180) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21322) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26573) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22967) * $signed(input_fmap_62[7:0]) +
	( 13'sd 4018) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28998) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21544) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_69[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7341) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27014) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8899) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11417) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26266) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5227) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21055) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20623) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17238) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11997) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30910) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20688) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2427) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10115) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18158) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16172) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14174) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26387) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25118) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2365) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21054) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1492) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7611) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22037) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11965) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20411) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11516) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22862) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11137) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25125) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_214;
assign conv_mac_214 = 
	( 15'sd 14537) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16128) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7812) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29432) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24284) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14045) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27046) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13729) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1885) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23994) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22987) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2765) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21654) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27233) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_16[7:0]) +
	( 10'sd 383) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6169) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7638) * $signed(input_fmap_21[7:0]) +
	( 10'sd 473) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12869) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5502) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31576) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27867) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32481) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2467) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16435) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13683) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15941) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24357) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29211) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29189) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13682) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2212) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28683) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21232) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10382) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29518) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4282) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5376) * $signed(input_fmap_51[7:0]) +
	( 8'sd 121) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19487) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23580) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32185) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8113) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1505) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30057) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24946) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20083) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15380) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16681) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20166) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23478) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17282) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9864) * $signed(input_fmap_70[7:0]) +
	( 9'sd 194) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16945) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16810) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28081) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6255) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9977) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4845) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10027) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31062) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24368) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15170) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30759) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24131) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18936) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27870) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21407) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1761) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12751) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16186) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29456) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23688) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26216) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31583) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12274) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29749) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1925) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20044) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5555) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21266) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17098) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7787) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4381) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12055) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31113) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27704) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9124) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24629) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2595) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16090) * $signed(input_fmap_123[7:0]) +
	( 14'sd 8112) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30656) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_215;
assign conv_mac_215 = 
	( 13'sd 3107) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25525) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3042) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30206) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22640) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7109) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8307) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19721) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32635) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16136) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7453) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9698) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5947) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7649) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15312) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10964) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9538) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28022) * $signed(input_fmap_28[7:0]) +
	( 11'sd 924) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29407) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31578) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29933) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17792) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2479) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19794) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13333) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12396) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4569) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1071) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32702) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6580) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2933) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16031) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24688) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28095) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11691) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5335) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5252) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27509) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31632) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1661) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22024) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30415) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20592) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1891) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14550) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10407) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29708) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21484) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_75[7:0]) +
	( 9'sd 232) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24620) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6965) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14300) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6663) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_82[7:0]) +
	( 9'sd 232) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11522) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3228) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15142) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28043) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28972) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15291) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24027) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15069) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21954) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11535) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4650) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10242) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24722) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16352) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18840) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19338) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4301) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20482) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3510) * $signed(input_fmap_107[7:0]) +
	( 7'sd 37) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22886) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20508) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23855) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19390) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12334) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14656) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8244) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8249) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27783) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20101) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_216;
assign conv_mac_216 = 
	( 13'sd 2187) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13019) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21732) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28024) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32138) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28594) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15015) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24274) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7923) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30427) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3873) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16383) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26736) * $signed(input_fmap_16[7:0]) +
	( 11'sd 582) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16853) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25651) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5281) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1357) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11411) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24206) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20364) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14156) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23786) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26323) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9700) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5051) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20055) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22260) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9275) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30381) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20505) * $signed(input_fmap_42[7:0]) +
	( 11'sd 781) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11950) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14486) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8504) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17415) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31057) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17372) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17884) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25979) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18936) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29667) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13318) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15011) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18302) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10630) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25534) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3287) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6887) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8390) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11592) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21962) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8899) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9214) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19575) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21492) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22398) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28865) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23692) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22795) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6309) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_83[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1081) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30790) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_87[7:0]) +
	( 9'sd 231) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14827) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11453) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22178) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27343) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1908) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19649) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24761) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30183) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22575) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31706) * $signed(input_fmap_102[7:0]) +
	( 11'sd 944) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7869) * $signed(input_fmap_104[7:0]) +
	( 11'sd 910) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22980) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17345) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32137) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28979) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6761) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3517) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18589) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29206) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26421) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8882) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23310) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17886) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27797) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24488) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_217;
assign conv_mac_217 = 
	( 16'sd 24618) * $signed(input_fmap_0[7:0]) +
	( 10'sd 501) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11520) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15826) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19976) * $signed(input_fmap_5[7:0]) +
	( 11'sd 567) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19386) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15389) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16617) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4727) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3337) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32281) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12063) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26025) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6079) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26809) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31079) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31990) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15440) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6880) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13020) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24165) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29644) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9740) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1610) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11080) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16181) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25371) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11863) * $signed(input_fmap_37[7:0]) +
	( 8'sd 121) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29533) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29089) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15402) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19005) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26562) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29350) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25397) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26731) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16830) * $signed(input_fmap_50[7:0]) +
	( 8'sd 101) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12609) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23578) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6730) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24110) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21663) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14197) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16873) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31851) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30522) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15971) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1859) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19794) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5456) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30204) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19049) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30457) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30900) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22961) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8816) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29350) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14819) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8178) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21187) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8540) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6739) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12893) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12393) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17859) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29522) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23785) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9290) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7608) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2739) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15791) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17744) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1110) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31192) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1028) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11475) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31111) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27068) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20202) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24975) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10742) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32165) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17665) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23046) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19854) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18486) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_218;
assign conv_mac_218 = 
	( 16'sd 18808) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12214) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30642) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28412) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10466) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27613) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27337) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26600) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25860) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13210) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22010) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8253) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14228) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_20[7:0]) +
	( 11'sd 886) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16218) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12835) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8618) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24765) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4360) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5947) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25736) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22602) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29520) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13913) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19288) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15405) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9198) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7157) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5905) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30969) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25935) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25839) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16827) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21228) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30255) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29831) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27678) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32492) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29290) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10042) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32451) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15727) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6589) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18743) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23684) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4439) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_70[7:0]) +
	( 10'sd 498) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29687) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5638) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28865) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28506) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28786) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27376) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21820) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9925) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12177) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31423) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22850) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21006) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10791) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25004) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7118) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13653) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30654) * $signed(input_fmap_98[7:0]) +
	( 12'sd 2001) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16338) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24073) * $signed(input_fmap_104[7:0]) +
	( 11'sd 537) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27529) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4456) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20971) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31458) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15931) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1039) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27408) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29312) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15353) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10973) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30596) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32664) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23544) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32193) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13313) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_219;
assign conv_mac_219 = 
	( 16'sd 28377) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25097) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12216) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5379) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29948) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3047) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2465) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9857) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6010) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28819) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25433) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30254) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19444) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11830) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5319) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26918) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31111) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22159) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27047) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32751) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13090) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4517) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8751) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26948) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16640) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13405) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23648) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21695) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7086) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3625) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14307) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25530) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1429) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21786) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15773) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6622) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9728) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19460) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30170) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11594) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15507) * $signed(input_fmap_73[7:0]) +
	( 14'sd 8048) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18382) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14201) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17442) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19729) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30206) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_85[7:0]) +
	( 10'sd 487) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22958) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11202) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2877) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16718) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23401) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19003) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30544) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29259) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10161) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30585) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27773) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32382) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1568) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12598) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20896) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20079) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12456) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26653) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5730) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2864) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21588) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24962) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3234) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7789) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_124[7:0]) +
	( 6'sd 23) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22114) * $signed(input_fmap_126[7:0]) +
	( 11'sd 558) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_220;
assign conv_mac_220 = 
	( 15'sd 15928) * $signed(input_fmap_0[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8888) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20946) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25276) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27339) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14639) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12052) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23891) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23076) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2559) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32019) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26552) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20996) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10501) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31601) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15548) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24911) * $signed(input_fmap_25[7:0]) +
	( 9'sd 220) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12355) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22736) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10432) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13236) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15156) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3367) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25439) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29066) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18029) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11851) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14699) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9350) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6114) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29275) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28551) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17446) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20823) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27680) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19721) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4877) * $signed(input_fmap_51[7:0]) +
	( 11'sd 906) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24195) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22057) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20919) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_61[7:0]) +
	( 7'sd 61) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21578) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19380) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29675) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30290) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7864) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32022) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13760) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13758) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26193) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28556) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20606) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21845) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6278) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8420) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1708) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18829) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18559) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21362) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2121) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19110) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9448) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8554) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17195) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4242) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25496) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19825) * $signed(input_fmap_110[7:0]) +
	( 11'sd 744) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13374) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32642) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31245) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32192) * $signed(input_fmap_116[7:0]) +
	( 5'sd 8) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22135) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_119[7:0]) +
	( 11'sd 794) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23017) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5845) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8277) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10747) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10009) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31455) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11151) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_221;
assign conv_mac_221 = 
	( 11'sd 630) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3205) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22087) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13581) * $signed(input_fmap_3[7:0]) +
	( 11'sd 642) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3479) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2868) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2633) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15321) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13414) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22069) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28221) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9931) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31403) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32619) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20631) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7647) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15488) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9170) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1571) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15987) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13351) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17157) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27285) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14634) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22925) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30332) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8733) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8776) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28024) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28005) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24746) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23061) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11888) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28942) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9240) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18431) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21561) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14582) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5030) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4416) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32537) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1147) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5134) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29921) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28131) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16280) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3631) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12124) * $signed(input_fmap_83[7:0]) +
	( 14'sd 8048) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14942) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25923) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27876) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3013) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20023) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28773) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4393) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4568) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32308) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29884) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1148) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16788) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15191) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6730) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12474) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14538) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15953) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6152) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27584) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8935) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28765) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2904) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22806) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13967) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14135) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27483) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4739) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25479) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_222;
assign conv_mac_222 = 
	( 15'sd 11455) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23257) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29024) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22856) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30394) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27507) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32658) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8155) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31900) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28266) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31739) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28448) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31935) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18564) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12200) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12460) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21885) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15656) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2054) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4779) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5855) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5926) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8028) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21995) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26308) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24156) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19369) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13170) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16356) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1085) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31271) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16645) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_49[7:0]) +
	( 11'sd 655) * $signed(input_fmap_50[7:0]) +
	( 10'sd 489) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11328) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22990) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24346) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6085) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9621) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7337) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12107) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11649) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3035) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27318) * $signed(input_fmap_62[7:0]) +
	( 9'sd 243) * $signed(input_fmap_63[7:0]) +
	( 10'sd 358) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16184) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_68[7:0]) +
	( 10'sd 269) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17722) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15453) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18688) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18522) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17445) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16355) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15036) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27684) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8964) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28502) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29852) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8412) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19590) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16942) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12161) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30272) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18256) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25068) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17003) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12110) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27472) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1884) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11633) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32201) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6547) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14112) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12461) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31198) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24321) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22702) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3126) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15596) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7014) * $signed(input_fmap_115[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10248) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19486) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26519) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27277) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3322) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6435) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_223;
assign conv_mac_223 = 
	( 15'sd 11615) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18687) * $signed(input_fmap_2[7:0]) +
	( 9'sd 207) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7436) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29117) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6970) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32005) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29346) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14791) * $signed(input_fmap_12[7:0]) +
	( 10'sd 269) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3593) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32476) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22885) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23854) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_20[7:0]) +
	( 13'sd 4009) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5827) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10605) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26647) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22968) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23110) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18368) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5819) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26662) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5999) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26705) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6496) * $signed(input_fmap_39[7:0]) +
	( 9'sd 245) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12157) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25122) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20060) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31303) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28204) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23699) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31892) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9738) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16143) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9368) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26373) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32028) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31545) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19749) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16581) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26904) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13784) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25537) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1090) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32443) * $signed(input_fmap_76[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27490) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14672) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30808) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31081) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15813) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9403) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17605) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8900) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7797) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29043) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20475) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7400) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9548) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28962) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13101) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5175) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22630) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15951) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12085) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23203) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9052) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31646) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5690) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27302) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10099) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32285) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19251) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15995) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_224;
assign conv_mac_224 = 
	( 16'sd 28066) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31513) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30811) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10213) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15517) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1970) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26024) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16576) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31461) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25345) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31465) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1809) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23399) * $signed(input_fmap_21[7:0]) +
	( 11'sd 591) * $signed(input_fmap_22[7:0]) +
	( 13'sd 4090) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21493) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23364) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17911) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22232) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14028) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20911) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16336) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26675) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25877) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18860) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26942) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27025) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7231) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24420) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18572) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18225) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2331) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29300) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19749) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16603) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22915) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28937) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1773) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16212) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6781) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2086) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17945) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26774) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27453) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29740) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31918) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17957) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16307) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2501) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4426) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4527) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20051) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1308) * $signed(input_fmap_78[7:0]) +
	( 11'sd 873) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29841) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26292) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30245) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19339) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19198) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7923) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24027) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3632) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23540) * $signed(input_fmap_97[7:0]) +
	( 9'sd 235) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11991) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26227) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29833) * $signed(input_fmap_101[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12185) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14740) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13939) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22026) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12071) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21238) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2819) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5551) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20653) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6387) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4975) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25700) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2892) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3021) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9454) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21159) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4387) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26601) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14027) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_225;
assign conv_mac_225 = 
	( 15'sd 14158) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17433) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6733) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31635) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14638) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27925) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18202) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11678) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15189) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11570) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6712) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17681) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5870) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7451) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2988) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24139) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12793) * $signed(input_fmap_23[7:0]) +
	( 9'sd 196) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29283) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13097) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16698) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19691) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18653) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2493) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18716) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26506) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24180) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14122) * $signed(input_fmap_39[7:0]) +
	( 11'sd 611) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6376) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29948) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26567) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27867) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9512) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8580) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18141) * $signed(input_fmap_49[7:0]) +
	( 9'sd 232) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19542) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30429) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9332) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18951) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24249) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20198) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23530) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16847) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26093) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24177) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25488) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6486) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14736) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11720) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16925) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22266) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19694) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5023) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7264) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3555) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_79[7:0]) +
	( 11'sd 684) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30049) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24714) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24287) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9471) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11779) * $signed(input_fmap_90[7:0]) +
	( 11'sd 990) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23674) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20800) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27450) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18680) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14642) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16361) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15015) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15710) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8275) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10396) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10691) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13548) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4785) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5156) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14845) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16953) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18725) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10033) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14950) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_116[7:0]) +
	( 11'sd 721) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23034) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30486) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27354) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14265) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4371) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30308) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_226;
assign conv_mac_226 = 
	( 10'sd 278) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10188) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25577) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1978) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4241) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11253) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24166) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_14[7:0]) +
	( 9'sd 130) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26164) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23048) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11395) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27167) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15375) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13447) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22413) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21087) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22335) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16233) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22353) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9490) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_35[7:0]) +
	( 10'sd 331) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29520) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28254) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1192) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16280) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19087) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8461) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11686) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30749) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32323) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2445) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15860) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13442) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1254) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12700) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19655) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8743) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15409) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12239) * $signed(input_fmap_65[7:0]) +
	( 8'sd 125) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9212) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9003) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22954) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17222) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8848) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31059) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18265) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6816) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21895) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27373) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18221) * $signed(input_fmap_86[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30577) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3263) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9809) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28522) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6326) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23852) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13532) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16433) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10747) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23668) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23821) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5231) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22372) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25348) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10460) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3484) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15488) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7626) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21221) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32035) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11312) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6072) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23331) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_227;
assign conv_mac_227 = 
	( 16'sd 16811) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23544) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8276) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9591) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7800) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6235) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29655) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12880) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1287) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11997) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24191) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30452) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28433) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31522) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24906) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24192) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23360) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4529) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16127) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30746) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22662) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7894) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8735) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26621) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6952) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15578) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30256) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1095) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9948) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23703) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9950) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10249) * $signed(input_fmap_48[7:0]) +
	( 12'sd 2008) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24637) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29004) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26034) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13688) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20900) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8544) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7078) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20783) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8806) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25274) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3298) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12593) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11319) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12722) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28039) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15029) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17966) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4719) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16762) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27475) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12288) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3419) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21390) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10390) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5942) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13591) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11306) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16500) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22788) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16999) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11584) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14830) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1059) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28577) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24856) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20247) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30100) * $signed(input_fmap_110[7:0]) +
	( 11'sd 591) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8725) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27908) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_115[7:0]) +
	( 8'sd 71) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19356) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13224) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19364) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_228;
assign conv_mac_228 = 
	( 15'sd 10994) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23804) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2543) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_3[7:0]) +
	( 13'sd 4075) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26564) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1604) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14625) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28686) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28213) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9420) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29746) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15222) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14606) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5901) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3921) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24423) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23854) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26907) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16477) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26013) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25057) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25567) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10029) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17807) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32675) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24461) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30202) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3264) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24716) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17839) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28559) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7991) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32001) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11265) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31278) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9998) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21424) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9311) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1313) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5141) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20482) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29503) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8820) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29850) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15015) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11031) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16556) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26929) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12665) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8318) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3631) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17252) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5667) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7880) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18126) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29689) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7914) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16203) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8301) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3667) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5024) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9783) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1796) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28618) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31319) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15103) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31822) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_94[7:0]) +
	( 11'sd 725) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25257) * $signed(input_fmap_96[7:0]) +
	( 11'sd 526) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26668) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5984) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17490) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8764) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6922) * $signed(input_fmap_104[7:0]) +
	( 9'sd 222) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10258) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19608) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18049) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_116[7:0]) +
	( 11'sd 977) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13516) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25322) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14790) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30504) * $signed(input_fmap_125[7:0]) +
	( 11'sd 619) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_229;
assign conv_mac_229 = 
	( 15'sd 12550) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14341) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7979) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13206) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25239) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1253) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12173) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26369) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24303) * $signed(input_fmap_19[7:0]) +
	( 14'sd 8165) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11855) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31221) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25921) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11252) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18121) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6124) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32040) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7362) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5176) * $signed(input_fmap_33[7:0]) +
	( 11'sd 691) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8254) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15212) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26004) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16809) * $signed(input_fmap_39[7:0]) +
	( 8'sd 103) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8266) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9609) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32537) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17664) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32349) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30089) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10545) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26741) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3289) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22913) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25972) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17331) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31083) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17969) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12985) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2577) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31005) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4142) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7517) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8348) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22600) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19000) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8619) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5895) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20086) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16798) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29180) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1145) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29409) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1152) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16418) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11072) * $signed(input_fmap_94[7:0]) +
	( 8'sd 83) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24201) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27297) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29265) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30405) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28201) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18142) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4309) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27985) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10728) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30426) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24072) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2490) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32251) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10395) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6405) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19952) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30346) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7725) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17769) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28366) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17998) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_230;
assign conv_mac_230 = 
	( 16'sd 31301) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25145) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6097) * $signed(input_fmap_3[7:0]) +
	( 10'sd 494) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10327) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16322) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10923) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8234) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18395) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25849) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27520) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31843) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27809) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3447) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28461) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27025) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6820) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10666) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3887) * $signed(input_fmap_29[7:0]) +
	( 11'sd 660) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11804) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5162) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4349) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1828) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1247) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23132) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_44[7:0]) +
	( 14'sd 8070) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22907) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6144) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23135) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30064) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12136) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25488) * $signed(input_fmap_52[7:0]) +
	( 11'sd 716) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21592) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5899) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21495) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7258) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23172) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5613) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10037) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4412) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2988) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21867) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23634) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13029) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12873) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11193) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19576) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22619) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19058) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17685) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27962) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23630) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31914) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22247) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17722) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11335) * $signed(input_fmap_88[7:0]) +
	( 10'sd 331) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4937) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26951) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9522) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12216) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22098) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6419) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17749) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31800) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18449) * $signed(input_fmap_101[7:0]) +
	( 12'sd 2005) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8723) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13964) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10397) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24646) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11028) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28241) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32400) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31770) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31573) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6989) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30296) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31887) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21957) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_231;
assign conv_mac_231 = 
	( 14'sd 4596) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6245) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17687) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8827) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17419) * $signed(input_fmap_5[7:0]) +
	( 9'sd 235) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32217) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12481) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29746) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12816) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23964) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31198) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3893) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28144) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23295) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20852) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15573) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9575) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18499) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13526) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5410) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6023) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19386) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7830) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30848) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3648) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18724) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27458) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20805) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8670) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23555) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17564) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3580) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30448) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5403) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28020) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4716) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9391) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7803) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14262) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18437) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1876) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16130) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19696) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9219) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28859) * $signed(input_fmap_71[7:0]) +
	( 10'sd 430) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29460) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29629) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32539) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9809) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18394) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17453) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18665) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27383) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3686) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27896) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24173) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14666) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11443) * $signed(input_fmap_93[7:0]) +
	( 14'sd 8123) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5383) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26922) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20562) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14861) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18475) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14675) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25617) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10464) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27912) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16662) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24202) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7626) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27190) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7752) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21877) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15708) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17624) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2762) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28197) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17378) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31693) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5742) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20601) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_232;
assign conv_mac_232 = 
	( 16'sd 28953) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20690) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16955) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1165) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5441) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6605) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11410) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1150) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14739) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17520) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29690) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11142) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9755) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19103) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32191) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11991) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1623) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17123) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1378) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31319) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2485) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10923) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28546) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24144) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19773) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29136) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27706) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18008) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4509) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15651) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14181) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3502) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32322) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19534) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15792) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5596) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29627) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3810) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10547) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28608) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2951) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16755) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28831) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23325) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4729) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19644) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16469) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2733) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17571) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24151) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5538) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14372) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4754) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31785) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7709) * $signed(input_fmap_90[7:0]) +
	( 10'sd 260) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8881) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28379) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17319) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26261) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9311) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8646) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_100[7:0]) +
	( 11'sd 831) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16489) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9706) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18043) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21169) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8456) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13788) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15866) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20682) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11793) * $signed(input_fmap_111[7:0]) +
	( 14'sd 8099) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5006) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21001) * $signed(input_fmap_115[7:0]) +
	( 11'sd 535) * $signed(input_fmap_116[7:0]) +
	( 11'sd 644) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17371) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7709) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21991) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25471) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21854) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14520) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4950) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_233;
assign conv_mac_233 = 
	( 16'sd 19735) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17272) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16971) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22790) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19537) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32520) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23126) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17474) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1258) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1410) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8926) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4980) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29938) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17965) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19690) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29277) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9261) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32073) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9783) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10237) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18482) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32180) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23418) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2383) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19530) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2663) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29922) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19073) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4918) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11320) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29124) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21965) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23555) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18660) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21175) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22819) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10198) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21880) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5622) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3479) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19015) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30154) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5603) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7584) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27948) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_75[7:0]) +
	( 11'sd 517) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16162) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_78[7:0]) +
	( 12'sd 2047) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1397) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18504) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7311) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10615) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1399) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14257) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12708) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3486) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26262) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29553) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4210) * $signed(input_fmap_97[7:0]) +
	( 12'sd 2039) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21860) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8444) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7982) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10541) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17677) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31608) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20307) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26034) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5762) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22983) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24401) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11577) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_115[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6067) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26651) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3828) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31741) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25685) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5879) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16052) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_234;
assign conv_mac_234 = 
	( 16'sd 29184) * $signed(input_fmap_0[7:0]) +
	( 10'sd 265) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27090) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22676) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18822) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12379) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28021) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11470) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18591) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28784) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16730) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4304) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11304) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21942) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20369) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9586) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11508) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24216) * $signed(input_fmap_28[7:0]) +
	( 10'sd 357) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5641) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29864) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17765) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24421) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13224) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3834) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11101) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_49[7:0]) +
	( 14'sd 8007) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12852) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3851) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32039) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5929) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6191) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32563) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2471) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3628) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17681) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30706) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8934) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10823) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7176) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2898) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14509) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27161) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30948) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32494) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22433) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_86[7:0]) +
	( 10'sd 420) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6242) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31954) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10128) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27132) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9871) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28200) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18635) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31275) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29555) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29349) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9240) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24299) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26188) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32455) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7007) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11438) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20927) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13376) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28904) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1872) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20703) * $signed(input_fmap_120[7:0]) +
	( 11'sd 590) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6530) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13752) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27839) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19436) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_235;
assign conv_mac_235 = 
	( 16'sd 19692) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20363) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1311) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28947) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2079) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31205) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18360) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_12[7:0]) +
	( 9'sd 150) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_14[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27213) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28681) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19081) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_20[7:0]) +
	( 11'sd 742) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1877) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28135) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24694) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21409) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6809) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11936) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1622) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7483) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_38[7:0]) +
	( 13'sd 4034) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17616) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4242) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2325) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5697) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19397) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22008) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26800) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28427) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16499) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2919) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7594) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11897) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1144) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18377) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7131) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24537) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1877) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6926) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14433) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16480) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4122) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28332) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_76[7:0]) +
	( 11'sd 983) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19407) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15254) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32026) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29801) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28181) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20426) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31286) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12789) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25074) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23439) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26677) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23539) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2121) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31783) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31629) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2396) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24397) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30251) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3872) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17385) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28960) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5124) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20025) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10587) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13243) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16543) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9435) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30344) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8127) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25286) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4444) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24410) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10057) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19040) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30337) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4590) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_236;
assign conv_mac_236 = 
	( 16'sd 29008) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13849) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28800) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4763) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17058) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22649) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24517) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26146) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16110) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17353) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21787) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6475) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3679) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20902) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3691) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28475) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20323) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7661) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6169) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27539) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32579) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1939) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26857) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27306) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1736) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12708) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25001) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16794) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20834) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10568) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4606) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11599) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21591) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31366) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22229) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5742) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23435) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17627) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5217) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18609) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13936) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28754) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3660) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21728) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21693) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19726) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18900) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18450) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23936) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29362) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31403) * $signed(input_fmap_97[7:0]) +
	( 6'sd 16) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4364) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27246) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28158) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9394) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7665) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28931) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20084) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26489) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1889) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31535) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12370) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3654) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30315) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32264) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14758) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8854) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22897) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31027) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30590) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23006) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32114) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7061) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_237;
assign conv_mac_237 = 
	( 16'sd 25289) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13259) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15519) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10338) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27907) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26049) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11652) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16827) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_17[7:0]) +
	( 11'sd 842) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32386) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23284) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8897) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31207) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24178) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25527) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31352) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30080) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15756) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30433) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30217) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25148) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22593) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6174) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14378) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7172) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14796) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10629) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32418) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26536) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31748) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16378) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8978) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_52[7:0]) +
	( 11'sd 987) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9948) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26582) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6995) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21362) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1148) * $signed(input_fmap_61[7:0]) +
	( 11'sd 690) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20099) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7630) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25049) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9937) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22679) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2218) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28789) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21840) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31347) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32075) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25669) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32179) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_77[7:0]) +
	( 10'sd 425) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27772) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29392) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11362) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21440) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29324) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23605) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27353) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14296) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12469) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28491) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6458) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5083) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10177) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8796) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27326) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9434) * $signed(input_fmap_110[7:0]) +
	( 9'sd 205) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13689) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9081) * $signed(input_fmap_114[7:0]) +
	( 11'sd 624) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8800) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6410) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22224) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5949) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3926) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30085) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2529) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23442) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_238;
assign conv_mac_238 = 
	( 16'sd 17077) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19027) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7694) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2053) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16926) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28269) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27691) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17424) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4862) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11237) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23149) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15620) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32081) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13173) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25206) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25858) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7296) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12552) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14919) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12448) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_37[7:0]) +
	( 11'sd 642) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32578) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24963) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18730) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18678) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29922) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30872) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28401) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13631) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11923) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24933) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15424) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2793) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14340) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31122) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32185) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24066) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2557) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_74[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17269) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11938) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16808) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16077) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9582) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21927) * $signed(input_fmap_84[7:0]) +
	( 11'sd 952) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24247) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11795) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22772) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3808) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12763) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4432) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32593) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6349) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28941) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7255) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13168) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9212) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22825) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18617) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4465) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14624) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1563) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27735) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17398) * $signed(input_fmap_110[7:0]) +
	( 11'sd 710) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19151) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8855) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23365) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3070) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24159) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11396) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8627) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28266) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9268) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_239;
assign conv_mac_239 = 
	( 16'sd 25851) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6573) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13490) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_4[7:0]) +
	( 11'sd 582) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21793) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15853) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4361) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20582) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9725) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8777) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29103) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9448) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30848) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9657) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2108) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10757) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18754) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30473) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23865) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27946) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10297) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5351) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11338) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3774) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19436) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22453) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14609) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25829) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25503) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30724) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5234) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_59[7:0]) +
	( 13'sd 4079) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24888) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21463) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13869) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9914) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27210) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19434) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14194) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14479) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12746) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11362) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11297) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27912) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11362) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25117) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23357) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20774) * $signed(input_fmap_85[7:0]) +
	( 9'sd 224) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15424) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9894) * $signed(input_fmap_89[7:0]) +
	( 8'sd 95) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21668) * $signed(input_fmap_91[7:0]) +
	( 8'sd 107) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13206) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11139) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23819) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7819) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12630) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5771) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31756) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8412) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4734) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7330) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22529) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11445) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13793) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27448) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12395) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14983) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12395) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32481) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13446) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24485) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_240;
assign conv_mac_240 = 
	( 14'sd 6058) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14147) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23287) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26601) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8299) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29255) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11589) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26898) * $signed(input_fmap_9[7:0]) +
	( 11'sd 540) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3246) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18118) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31818) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3854) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30594) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2297) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25472) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2160) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16158) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1813) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28910) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10884) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17669) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12597) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21999) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24467) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7761) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21455) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3783) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27199) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4953) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21306) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3962) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20323) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26262) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17120) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7679) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19909) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16050) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6892) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18163) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32516) * $signed(input_fmap_53[7:0]) +
	( 11'sd 807) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24998) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8477) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16149) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7336) * $signed(input_fmap_59[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19607) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2398) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15039) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17328) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25526) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14256) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14831) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29705) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5584) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11448) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17982) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20374) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18402) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15202) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25947) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25387) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3152) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14218) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29202) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7238) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23185) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4643) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26838) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12344) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_96[7:0]) +
	( 11'sd 555) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20843) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13202) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18661) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12839) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11231) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21520) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31911) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10219) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19619) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9628) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22899) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19295) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11760) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_120[7:0]) +
	( 11'sd 869) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15501) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2699) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2065) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12809) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_241;
assign conv_mac_241 = 
	( 16'sd 16518) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26453) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7285) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11102) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30536) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3417) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23694) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14910) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1817) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12404) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30328) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25624) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26916) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13804) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29487) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30625) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21903) * $signed(input_fmap_33[7:0]) +
	( 10'sd 382) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10046) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5745) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5217) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2935) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23601) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21966) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14269) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28654) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30558) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20794) * $signed(input_fmap_46[7:0]) +
	( 12'sd 2030) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6351) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26198) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31374) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30705) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28622) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29043) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22564) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2649) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18975) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4128) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23546) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29306) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6932) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13906) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25188) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30119) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22338) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23653) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6611) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17857) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13453) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10376) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15781) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21837) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16609) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17606) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2396) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28048) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11457) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29356) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19385) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12331) * $signed(input_fmap_104[7:0]) +
	( 11'sd 731) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17700) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18256) * $signed(input_fmap_108[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16879) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9154) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17277) * $signed(input_fmap_113[7:0]) +
	( 10'sd 438) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2832) * $signed(input_fmap_115[7:0]) +
	( 11'sd 616) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17180) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12062) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3489) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9548) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16014) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19892) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14940) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_242;
assign conv_mac_242 = 
	( 13'sd 3188) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27470) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30601) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21277) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5158) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3350) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30811) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9765) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5634) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15396) * $signed(input_fmap_16[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8783) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14910) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16251) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12221) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2303) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25313) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6581) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20742) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6467) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14074) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14578) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13315) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4515) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2691) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28427) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32167) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19589) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12936) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6249) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2514) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1888) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2482) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12032) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12396) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28745) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23639) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19740) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24261) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11398) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16476) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23746) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13166) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6213) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27407) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9249) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3179) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24757) * $signed(input_fmap_70[7:0]) +
	( 8'sd 118) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21017) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26414) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_78[7:0]) +
	( 9'sd 183) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26034) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32291) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27884) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21772) * $signed(input_fmap_86[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1410) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6395) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9183) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1477) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17360) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_98[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4113) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4687) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10876) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21551) * $signed(input_fmap_107[7:0]) +
	( 5'sd 12) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27723) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32586) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_112[7:0]) +
	( 9'sd 203) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7307) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13408) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9553) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13023) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31600) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26373) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_243;
assign conv_mac_243 = 
	( 16'sd 25018) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30345) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27882) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29017) * $signed(input_fmap_4[7:0]) +
	( 11'sd 619) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18390) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15762) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32755) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23446) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28621) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17786) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8939) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3824) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16487) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4238) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1227) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30890) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10053) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13942) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29116) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2617) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19821) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24723) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28006) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25458) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28394) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22042) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24369) * $signed(input_fmap_37[7:0]) +
	( 11'sd 722) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15425) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15459) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22763) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28875) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26656) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1338) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11563) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12801) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13696) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28410) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9420) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11036) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10776) * $signed(input_fmap_55[7:0]) +
	( 11'sd 545) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21472) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7733) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23734) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6182) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22550) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30074) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_66[7:0]) +
	( 13'sd 4002) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24802) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18896) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25257) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26901) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19247) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29938) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32021) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30198) * $signed(input_fmap_77[7:0]) +
	( 11'sd 782) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24262) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2441) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15194) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29776) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5132) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7100) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2128) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5995) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1938) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7730) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6675) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13181) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7168) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4834) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25027) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12942) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32497) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15235) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6943) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9098) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23793) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30193) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6859) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7115) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26375) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16958) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13199) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13127) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32117) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32546) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28347) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_244;
assign conv_mac_244 = 
	( 16'sd 25461) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10593) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25860) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9038) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22307) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24303) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10630) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26587) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2683) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14091) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6855) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10732) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3305) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3253) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20411) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13478) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16619) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23349) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10635) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16313) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19267) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23390) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27399) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31717) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3339) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3045) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28294) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20277) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7422) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6727) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9825) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24995) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8875) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14237) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9595) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14925) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10647) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9105) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18064) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6025) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26813) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17374) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13437) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27578) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23645) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24197) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14024) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27400) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23626) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20183) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12708) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_88[7:0]) +
	( 6'sd 31) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3274) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3310) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25749) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19973) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6383) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14561) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5155) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29184) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28773) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_100[7:0]) +
	( 8'sd 71) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26968) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18347) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22017) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13236) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23315) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19224) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27608) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21464) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14658) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11053) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11774) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7274) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9256) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31626) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13102) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18766) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9085) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29417) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26028) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_245;
assign conv_mac_245 = 
	( 16'sd 23574) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25968) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11261) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11231) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5720) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_8[7:0]) +
	( 13'sd 4046) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22816) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30225) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6152) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15648) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31875) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1313) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23541) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1811) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16768) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2451) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5180) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18635) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26841) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5223) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15295) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12988) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15079) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13316) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26113) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18706) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11890) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_46[7:0]) +
	( 11'sd 586) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24824) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11797) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24156) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19197) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13148) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12378) * $signed(input_fmap_63[7:0]) +
	( 11'sd 577) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13458) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15819) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10955) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24067) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21292) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29015) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11515) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25519) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6186) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4623) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15010) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18769) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25083) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24067) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9721) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29068) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25340) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30727) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4722) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31493) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3469) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29011) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2852) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26307) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16712) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4898) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24598) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28371) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2371) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32547) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16375) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32060) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7080) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10339) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_115[7:0]) +
	( 10'sd 378) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24602) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27908) * $signed(input_fmap_120[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8779) * $signed(input_fmap_122[7:0]) +
	( 8'sd 90) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7095) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23756) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7167) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14172) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_246;
assign conv_mac_246 = 
	( 16'sd 18001) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20277) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9661) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12770) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1119) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24793) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5772) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24400) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12042) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10411) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1888) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22530) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20504) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26882) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18262) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26376) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26805) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19362) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20714) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21505) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24032) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23032) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_29[7:0]) +
	( 11'sd 826) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31457) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22437) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27285) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28760) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18183) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23429) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5585) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23911) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10964) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16206) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9687) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23288) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16541) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26290) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19462) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16055) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_62[7:0]) +
	( 10'sd 315) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7916) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24201) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4207) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27425) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26226) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22542) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27935) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27207) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29287) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3787) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20996) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20878) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17277) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23013) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29633) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19236) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22468) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10436) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14136) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25125) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5945) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9846) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5431) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14145) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21980) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2692) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25408) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8508) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23153) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30414) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7875) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24749) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_122[7:0]) +
	( 7'sd 56) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24271) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_247;
assign conv_mac_247 = 
	( 11'sd 927) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14321) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11938) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23067) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29203) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3795) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14167) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24593) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29031) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15720) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11607) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19826) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28550) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23371) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2108) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8453) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28974) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28876) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17606) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21298) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12060) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29522) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7542) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26770) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24610) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31348) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21807) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2118) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29502) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14085) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24027) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9341) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13705) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22956) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26831) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28711) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28596) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30857) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23355) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11364) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15939) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7155) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5352) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22158) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3217) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25680) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_67[7:0]) +
	( 10'sd 324) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3986) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17465) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4449) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15167) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10301) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19103) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24902) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29224) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25233) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27638) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15566) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25802) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10972) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16910) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8238) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8512) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27600) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1477) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32056) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17248) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2050) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21993) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1083) * $signed(input_fmap_103[7:0]) +
	( 11'sd 1022) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30146) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19914) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27014) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32301) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18300) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15289) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23622) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6799) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24782) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15204) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24642) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12034) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4267) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22382) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4953) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3322) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17561) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14478) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_248;
assign conv_mac_248 = 
	( 13'sd 3905) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23272) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4404) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20933) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29863) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16753) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6499) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1259) * $signed(input_fmap_11[7:0]) +
	( 11'sd 550) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31865) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16241) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27671) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4959) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1349) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16148) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11972) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_24[7:0]) +
	( 10'sd 473) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23729) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13977) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4327) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26367) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29041) * $signed(input_fmap_31[7:0]) +
	( 11'sd 859) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1657) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3356) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17744) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30077) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24016) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16105) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15609) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10792) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6376) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7176) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27723) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31303) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23463) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16844) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18669) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29136) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22285) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29825) * $signed(input_fmap_57[7:0]) +
	( 11'sd 962) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8472) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26549) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19972) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5500) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18770) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6355) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27212) * $signed(input_fmap_68[7:0]) +
	( 10'sd 354) * $signed(input_fmap_69[7:0]) +
	( 10'sd 343) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10941) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12423) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14053) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1365) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2697) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4416) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14078) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1195) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22988) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8524) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27338) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27252) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15301) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25094) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5202) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_96[7:0]) +
	( 9'sd 192) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31211) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15255) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29865) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20303) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6154) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10078) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7089) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29979) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22237) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25450) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9938) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13801) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1240) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8313) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3529) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7328) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10691) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31362) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21921) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_249;
assign conv_mac_249 = 
	( 15'sd 14011) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_1[7:0]) +
	( 11'sd 691) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20973) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19867) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32440) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3096) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31078) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13122) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22184) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27699) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28677) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31105) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2308) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13391) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28023) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21706) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30506) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_26[7:0]) +
	( 11'sd 984) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21066) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11756) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11368) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13505) * $signed(input_fmap_33[7:0]) +
	( 10'sd 305) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23952) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2924) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23002) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32482) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26746) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15948) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4881) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4143) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12854) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28393) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5896) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28273) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29051) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16860) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28675) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23370) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21480) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7829) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15062) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30820) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22308) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24299) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3348) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31237) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1723) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32141) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31500) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18409) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21993) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7820) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2899) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12615) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15610) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11951) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15824) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32243) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30078) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19812) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5463) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22074) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10595) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4480) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1140) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19302) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3361) * $signed(input_fmap_102[7:0]) +
	( 11'sd 724) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19005) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10872) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3467) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15227) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18080) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9831) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2475) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13184) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12481) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8023) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22819) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23316) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6100) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25910) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22875) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30261) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13538) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14547) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_250;
assign conv_mac_250 = 
	( 15'sd 8878) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30927) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15478) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26180) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13738) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10875) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23386) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15399) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24776) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19984) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25715) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19699) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25942) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25851) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19542) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2300) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31535) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9378) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9738) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26634) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11766) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32026) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30235) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6214) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17310) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2455) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32068) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12539) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4711) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20239) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4961) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20969) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15144) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3620) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18282) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12984) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10451) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15079) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_56[7:0]) +
	( 11'sd 908) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9381) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10345) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3600) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1099) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2355) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11319) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13532) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21657) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11484) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7658) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30261) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26076) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15925) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14781) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20726) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8443) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31571) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26566) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7761) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24041) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30736) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19219) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10784) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14942) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6306) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10860) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7461) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18154) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9478) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14500) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31954) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2054) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27675) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15538) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32397) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28470) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14205) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22803) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11071) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8429) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27774) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7276) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23403) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8634) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15155) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_251;
assign conv_mac_251 = 
	( 16'sd 30875) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16486) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6367) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8638) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13271) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14059) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6933) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3671) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17790) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13061) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16989) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28577) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32694) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23593) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10307) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2994) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6306) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1726) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25170) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13110) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8828) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25657) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5169) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3230) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21789) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30783) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20190) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_44[7:0]) +
	( 11'sd 599) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14838) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29722) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7322) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31782) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3684) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1671) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_54[7:0]) +
	( 11'sd 854) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23713) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25170) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18256) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14065) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5086) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13247) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27220) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9937) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11519) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24306) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15759) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8607) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31071) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28141) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26470) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29624) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17835) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31812) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4742) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21034) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1947) * $signed(input_fmap_85[7:0]) +
	( 8'sd 102) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32701) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28331) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10585) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6762) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10644) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14504) * $signed(input_fmap_93[7:0]) +
	( 11'sd 608) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13418) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24156) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2642) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14882) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18570) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27231) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28539) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25906) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5057) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27222) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21452) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18453) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15765) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1189) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1675) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31746) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17055) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2994) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30548) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_252;
assign conv_mac_252 = 
	( 15'sd 9572) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26018) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23131) * $signed(input_fmap_2[7:0]) +
	( 11'sd 602) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9899) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24614) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30753) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7195) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25357) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24658) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27259) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3619) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3444) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27477) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20730) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30346) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28540) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3061) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16440) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9473) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25665) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7177) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12972) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11901) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11498) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19428) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21763) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16761) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8807) * $signed(input_fmap_48[7:0]) +
	( 11'sd 952) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24225) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2393) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25433) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16573) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11801) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12444) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31051) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12673) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27774) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21185) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3350) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10998) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6627) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3619) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27576) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18599) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24523) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3034) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13003) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19379) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16182) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29514) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9573) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22080) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28514) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14402) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11434) * $signed(input_fmap_97[7:0]) +
	( 11'sd 613) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10129) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10082) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16083) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11853) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27662) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25952) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29814) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24711) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2921) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7066) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29278) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11984) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25620) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21353) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31995) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29994) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28867) * $signed(input_fmap_126[7:0]) +
	( 7'sd 54) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_253;
assign conv_mac_253 = 
	( 16'sd 24828) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24192) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30969) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4656) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10005) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14351) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24644) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11770) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26842) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6686) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5235) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14942) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32054) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27937) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28765) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30509) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32484) * $signed(input_fmap_19[7:0]) +
	( 9'sd 198) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8607) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26324) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10668) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9610) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1573) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19028) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21078) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16092) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17802) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8042) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17239) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17747) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9526) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28271) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16602) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19033) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23141) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15901) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3512) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25791) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7888) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30456) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3298) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20006) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19307) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23951) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23665) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26745) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26375) * $signed(input_fmap_62[7:0]) +
	( 11'sd 939) * $signed(input_fmap_63[7:0]) +
	( 9'sd 161) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25215) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8179) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3242) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22990) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26124) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2283) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3144) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20381) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23988) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30725) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20354) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15768) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21682) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23788) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12811) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30404) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25475) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20505) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30391) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2419) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5786) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_92[7:0]) +
	( 11'sd 793) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10153) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31655) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14999) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30619) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18147) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5443) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20566) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14826) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13269) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1951) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8239) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9776) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22485) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26189) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16358) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16214) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18383) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26895) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_119[7:0]) +
	( 10'sd 493) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8489) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20764) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17182) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26557) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_254;
assign conv_mac_254 = 
	( 15'sd 8728) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27983) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30688) * $signed(input_fmap_2[7:0]) +
	( 9'sd 241) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9334) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5344) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24681) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27609) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_10[7:0]) +
	( 11'sd 611) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13647) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21888) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31226) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5048) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32723) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11420) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20194) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9448) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25171) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12257) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4152) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6429) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11570) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18960) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13885) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13730) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21066) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_44[7:0]) +
	( 9'sd 252) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13817) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14280) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7325) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21805) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30642) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30106) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9248) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26353) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14538) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12980) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31224) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2684) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19272) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18875) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12508) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3709) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8523) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19888) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30033) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6542) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8941) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13227) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23330) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4475) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11111) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19170) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1414) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9976) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23157) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22846) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8847) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2691) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26567) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12256) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19395) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21256) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1813) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_103[7:0]) +
	( 10'sd 352) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12601) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2255) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7908) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18785) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16836) * $signed(input_fmap_110[7:0]) +
	( 10'sd 256) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31470) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21700) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1097) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10873) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12525) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25241) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23581) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13401) * $signed(input_fmap_120[7:0]) +
	( 9'sd 186) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19665) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12372) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4778) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11300) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_255;
assign conv_mac_255 = 
	( 16'sd 29970) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11486) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22690) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11542) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20368) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10660) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3641) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24756) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4813) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30575) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12071) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2783) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1283) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27648) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31594) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13414) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_24[7:0]) +
	( 9'sd 185) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23162) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24054) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20047) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10795) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17675) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25729) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2880) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9368) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28501) * $signed(input_fmap_37[7:0]) +
	( 10'sd 505) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27569) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7662) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31075) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26966) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2907) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8459) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17779) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10421) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6786) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15962) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14084) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2704) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27562) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28180) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4263) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25260) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23695) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20180) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12293) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3897) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5195) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12751) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32588) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13157) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13007) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19064) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30279) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25473) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7269) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4516) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4585) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20165) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6194) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19213) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16377) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2766) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10756) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1562) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23923) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22509) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32012) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14464) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5109) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_111[7:0]) +
	( 14'sd 8186) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14298) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4586) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16447) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5311) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24504) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23708) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6005) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5230) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29127) * $signed(input_fmap_127[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 16'd20546;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 16'd20498;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 15'd13188;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 15'd16181;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 15'd14581;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 16'd21931;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 16'd22488;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 11'd561;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 15'd11003;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 16'd24987;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 16'd23492;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 16'd19197;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 15'd8619;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 14'd4771;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 16'd24075;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 16'd18603;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 15'd15259;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 16'd31604;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 14'd6815;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 16'd18522;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 15'd8610;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 14'd5435;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 15'd10250;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 16'd21566;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 15'd14283;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 14'd6995;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 16'd28747;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 11'd724;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 16'd28522;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 14'd5560;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 14'd4668;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 15'd9754;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 15'd12389;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 16'd21626;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 12'd1346;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 16'd20698;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 16'd19256;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 14'd8103;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 15'd16000;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 16'd19714;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 16'd16920;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 14'd4254;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 16'd29005;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 15'd9698;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 14'd6668;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 11'd630;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 15'd12641;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 10'd278;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 13'd3352;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 16'd18686;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 14'd4845;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 15'd11086;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 15'd11543;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 16'd28314;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 16'd18116;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 16'd30260;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 14'd5793;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 16'd29254;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 15'd9126;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 9'd166;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 15'd10149;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 16'd24001;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 15'd10443;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 16'd24051;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 13'd3445;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 15'd8926;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 15'd16376;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 13'd3095;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 16'd22860;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 15'd13187;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 15'd8644;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 11'd964;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 16'd23445;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 15'd9454;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 16'd29390;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 11'd758;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 15'd8416;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 15'd13048;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 11'd807;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 14'd8035;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 14'd4757;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 16'd26146;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 16'd26078;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 15'd10114;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 16'd32481;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 13'd2539;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 15'd9327;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 16'd19078;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 16'd20324;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 15'd9159;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 15'd13263;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 16'd28740;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 15'd8885;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 16'd28080;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 16'd32198;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 16'd31428;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 16'd28126;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 14'd4788;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 16'd32357;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 16'd29690;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 12'd1586;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 16'd28716;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 16'd16437;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 16'd28449;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 16'd32014;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 16'd26912;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 16'd23864;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 16'd23156;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 13'd2419;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 15'd9708;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 16'd22070;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 16'd21042;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 15'd13303;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 16'd19568;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 13'd3037;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 15'd12110;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 15'd13529;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 16'd25005;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 16'd17249;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 14'd4317;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 16'd23881;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 15'd9795;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 16'd18202;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 15'd12905;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 14'd5570;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 14'd4099;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 16'd28048;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 16'd31743;
logic [31:0] bias_add_128;
assign bias_add_128 = conv_mac_128 + 15'd12348;
logic [31:0] bias_add_129;
assign bias_add_129 = conv_mac_129 + 16'd18592;
logic [31:0] bias_add_130;
assign bias_add_130 = conv_mac_130 + 16'd28157;
logic [31:0] bias_add_131;
assign bias_add_131 = conv_mac_131 + 16'd32347;
logic [31:0] bias_add_132;
assign bias_add_132 = conv_mac_132 + 16'd16397;
logic [31:0] bias_add_133;
assign bias_add_133 = conv_mac_133 + 12'd1148;
logic [31:0] bias_add_134;
assign bias_add_134 = conv_mac_134 + 15'd12203;
logic [31:0] bias_add_135;
assign bias_add_135 = conv_mac_135 + 16'd25952;
logic [31:0] bias_add_136;
assign bias_add_136 = conv_mac_136 + 16'd31141;
logic [31:0] bias_add_137;
assign bias_add_137 = conv_mac_137 + 14'd5651;
logic [31:0] bias_add_138;
assign bias_add_138 = conv_mac_138 + 16'd18145;
logic [31:0] bias_add_139;
assign bias_add_139 = conv_mac_139 + 14'd5086;
logic [31:0] bias_add_140;
assign bias_add_140 = conv_mac_140 + 16'd18153;
logic [31:0] bias_add_141;
assign bias_add_141 = conv_mac_141 + 16'd20847;
logic [31:0] bias_add_142;
assign bias_add_142 = conv_mac_142 + 15'd15109;
logic [31:0] bias_add_143;
assign bias_add_143 = conv_mac_143 + 15'd16005;
logic [31:0] bias_add_144;
assign bias_add_144 = conv_mac_144 + 15'd12978;
logic [31:0] bias_add_145;
assign bias_add_145 = conv_mac_145 + 14'd7990;
logic [31:0] bias_add_146;
assign bias_add_146 = conv_mac_146 + 13'd3266;
logic [31:0] bias_add_147;
assign bias_add_147 = conv_mac_147 + 16'd25077;
logic [31:0] bias_add_148;
assign bias_add_148 = conv_mac_148 + 16'd26644;
logic [31:0] bias_add_149;
assign bias_add_149 = conv_mac_149 + 15'd14683;
logic [31:0] bias_add_150;
assign bias_add_150 = conv_mac_150 + 15'd8854;
logic [31:0] bias_add_151;
assign bias_add_151 = conv_mac_151 + 16'd22890;
logic [31:0] bias_add_152;
assign bias_add_152 = conv_mac_152 + 16'd27105;
logic [31:0] bias_add_153;
assign bias_add_153 = conv_mac_153 + 15'd11302;
logic [31:0] bias_add_154;
assign bias_add_154 = conv_mac_154 + 15'd13185;
logic [31:0] bias_add_155;
assign bias_add_155 = conv_mac_155 + 16'd27242;
logic [31:0] bias_add_156;
assign bias_add_156 = conv_mac_156 + 15'd8457;
logic [31:0] bias_add_157;
assign bias_add_157 = conv_mac_157 + 16'd19223;
logic [31:0] bias_add_158;
assign bias_add_158 = conv_mac_158 + 15'd15884;
logic [31:0] bias_add_159;
assign bias_add_159 = conv_mac_159 + 14'd7316;
logic [31:0] bias_add_160;
assign bias_add_160 = conv_mac_160 + 16'd22042;
logic [31:0] bias_add_161;
assign bias_add_161 = conv_mac_161 + 13'd3803;
logic [31:0] bias_add_162;
assign bias_add_162 = conv_mac_162 + 16'd26258;
logic [31:0] bias_add_163;
assign bias_add_163 = conv_mac_163 + 13'd2473;
logic [31:0] bias_add_164;
assign bias_add_164 = conv_mac_164 + 14'd4155;
logic [31:0] bias_add_165;
assign bias_add_165 = conv_mac_165 + 16'd20443;
logic [31:0] bias_add_166;
assign bias_add_166 = conv_mac_166 + 10'd334;
logic [31:0] bias_add_167;
assign bias_add_167 = conv_mac_167 + 16'd17036;
logic [31:0] bias_add_168;
assign bias_add_168 = conv_mac_168 + 12'd1593;
logic [31:0] bias_add_169;
assign bias_add_169 = conv_mac_169 + 15'd15000;
logic [31:0] bias_add_170;
assign bias_add_170 = conv_mac_170 + 14'd4708;
logic [31:0] bias_add_171;
assign bias_add_171 = conv_mac_171 + 15'd9663;
logic [31:0] bias_add_172;
assign bias_add_172 = conv_mac_172 + 14'd5709;
logic [31:0] bias_add_173;
assign bias_add_173 = conv_mac_173 + 16'd29889;
logic [31:0] bias_add_174;
assign bias_add_174 = conv_mac_174 + 14'd6415;
logic [31:0] bias_add_175;
assign bias_add_175 = conv_mac_175 + 16'd29068;
logic [31:0] bias_add_176;
assign bias_add_176 = conv_mac_176 + 16'd21017;
logic [31:0] bias_add_177;
assign bias_add_177 = conv_mac_177 + 14'd4667;
logic [31:0] bias_add_178;
assign bias_add_178 = conv_mac_178 + 14'd6005;
logic [31:0] bias_add_179;
assign bias_add_179 = conv_mac_179 + 16'd26955;
logic [31:0] bias_add_180;
assign bias_add_180 = conv_mac_180 + 12'd1403;
logic [31:0] bias_add_181;
assign bias_add_181 = conv_mac_181 + 13'd2818;
logic [31:0] bias_add_182;
assign bias_add_182 = conv_mac_182 + 16'd24924;
logic [31:0] bias_add_183;
assign bias_add_183 = conv_mac_183 + 14'd5787;
logic [31:0] bias_add_184;
assign bias_add_184 = conv_mac_184 + 15'd9555;
logic [31:0] bias_add_185;
assign bias_add_185 = conv_mac_185 + 16'd18155;
logic [31:0] bias_add_186;
assign bias_add_186 = conv_mac_186 + 12'd1743;
logic [31:0] bias_add_187;
assign bias_add_187 = conv_mac_187 + 16'd21530;
logic [31:0] bias_add_188;
assign bias_add_188 = conv_mac_188 + 16'd27847;
logic [31:0] bias_add_189;
assign bias_add_189 = conv_mac_189 + 16'd22850;
logic [31:0] bias_add_190;
assign bias_add_190 = conv_mac_190 + 16'd29355;
logic [31:0] bias_add_191;
assign bias_add_191 = conv_mac_191 + 13'd2606;
logic [31:0] bias_add_192;
assign bias_add_192 = conv_mac_192 + 16'd20677;
logic [31:0] bias_add_193;
assign bias_add_193 = conv_mac_193 + 12'd1993;
logic [31:0] bias_add_194;
assign bias_add_194 = conv_mac_194 + 12'd1680;
logic [31:0] bias_add_195;
assign bias_add_195 = conv_mac_195 + 16'd30259;
logic [31:0] bias_add_196;
assign bias_add_196 = conv_mac_196 + 16'd27720;
logic [31:0] bias_add_197;
assign bias_add_197 = conv_mac_197 + 15'd8207;
logic [31:0] bias_add_198;
assign bias_add_198 = conv_mac_198 + 15'd11283;
logic [31:0] bias_add_199;
assign bias_add_199 = conv_mac_199 + 14'd8129;
logic [31:0] bias_add_200;
assign bias_add_200 = conv_mac_200 + 16'd31305;
logic [31:0] bias_add_201;
assign bias_add_201 = conv_mac_201 + 14'd8170;
logic [31:0] bias_add_202;
assign bias_add_202 = conv_mac_202 + 14'd6397;
logic [31:0] bias_add_203;
assign bias_add_203 = conv_mac_203 + 15'd15540;
logic [31:0] bias_add_204;
assign bias_add_204 = conv_mac_204 + 16'd18240;
logic [31:0] bias_add_205;
assign bias_add_205 = conv_mac_205 + 15'd15046;
logic [31:0] bias_add_206;
assign bias_add_206 = conv_mac_206 + 16'd23646;
logic [31:0] bias_add_207;
assign bias_add_207 = conv_mac_207 + 13'd3612;
logic [31:0] bias_add_208;
assign bias_add_208 = conv_mac_208 + 16'd22303;
logic [31:0] bias_add_209;
assign bias_add_209 = conv_mac_209 + 14'd5228;
logic [31:0] bias_add_210;
assign bias_add_210 = conv_mac_210 + 15'd11261;
logic [31:0] bias_add_211;
assign bias_add_211 = conv_mac_211 + 16'd19876;
logic [31:0] bias_add_212;
assign bias_add_212 = conv_mac_212 + 15'd15835;
logic [31:0] bias_add_213;
assign bias_add_213 = conv_mac_213 + 16'd29397;
logic [31:0] bias_add_214;
assign bias_add_214 = conv_mac_214 + 15'd13577;
logic [31:0] bias_add_215;
assign bias_add_215 = conv_mac_215 + 15'd14402;
logic [31:0] bias_add_216;
assign bias_add_216 = conv_mac_216 + 15'd11424;
logic [31:0] bias_add_217;
assign bias_add_217 = conv_mac_217 + 11'd801;
logic [31:0] bias_add_218;
assign bias_add_218 = conv_mac_218 + 15'd16046;
logic [31:0] bias_add_219;
assign bias_add_219 = conv_mac_219 + 16'd31640;
logic [31:0] bias_add_220;
assign bias_add_220 = conv_mac_220 + 15'd11406;
logic [31:0] bias_add_221;
assign bias_add_221 = conv_mac_221 + 16'd23359;
logic [31:0] bias_add_222;
assign bias_add_222 = conv_mac_222 + 16'd32028;
logic [31:0] bias_add_223;
assign bias_add_223 = conv_mac_223 + 12'd1818;
logic [31:0] bias_add_224;
assign bias_add_224 = conv_mac_224 + 15'd12452;
logic [31:0] bias_add_225;
assign bias_add_225 = conv_mac_225 + 16'd20922;
logic [31:0] bias_add_226;
assign bias_add_226 = conv_mac_226 + 16'd20603;
logic [31:0] bias_add_227;
assign bias_add_227 = conv_mac_227 + 15'd8323;
logic [31:0] bias_add_228;
assign bias_add_228 = conv_mac_228 + 15'd13400;
logic [31:0] bias_add_229;
assign bias_add_229 = conv_mac_229 + 15'd10299;
logic [31:0] bias_add_230;
assign bias_add_230 = conv_mac_230 + 13'd2458;
logic [31:0] bias_add_231;
assign bias_add_231 = conv_mac_231 + 13'd3523;
logic [31:0] bias_add_232;
assign bias_add_232 = conv_mac_232 + 16'd25672;
logic [31:0] bias_add_233;
assign bias_add_233 = conv_mac_233 + 16'd26104;
logic [31:0] bias_add_234;
assign bias_add_234 = conv_mac_234 + 16'd20355;
logic [31:0] bias_add_235;
assign bias_add_235 = conv_mac_235 + 16'd19505;
logic [31:0] bias_add_236;
assign bias_add_236 = conv_mac_236 + 16'd31731;
logic [31:0] bias_add_237;
assign bias_add_237 = conv_mac_237 + 16'd29947;
logic [31:0] bias_add_238;
assign bias_add_238 = conv_mac_238 + 16'd29142;
logic [31:0] bias_add_239;
assign bias_add_239 = conv_mac_239 + 15'd13778;
logic [31:0] bias_add_240;
assign bias_add_240 = conv_mac_240 + 7'd39;
logic [31:0] bias_add_241;
assign bias_add_241 = conv_mac_241 + 16'd21171;
logic [31:0] bias_add_242;
assign bias_add_242 = conv_mac_242 + 16'd19039;
logic [31:0] bias_add_243;
assign bias_add_243 = conv_mac_243 + 16'd17452;
logic [31:0] bias_add_244;
assign bias_add_244 = conv_mac_244 + 16'd20322;
logic [31:0] bias_add_245;
assign bias_add_245 = conv_mac_245 + 16'd21028;
logic [31:0] bias_add_246;
assign bias_add_246 = conv_mac_246 + 15'd10934;
logic [31:0] bias_add_247;
assign bias_add_247 = conv_mac_247 + 16'd21564;
logic [31:0] bias_add_248;
assign bias_add_248 = conv_mac_248 + 16'd20133;
logic [31:0] bias_add_249;
assign bias_add_249 = conv_mac_249 + 15'd9249;
logic [31:0] bias_add_250;
assign bias_add_250 = conv_mac_250 + 16'd17198;
logic [31:0] bias_add_251;
assign bias_add_251 = conv_mac_251 + 15'd10231;
logic [31:0] bias_add_252;
assign bias_add_252 = conv_mac_252 + 16'd17284;
logic [31:0] bias_add_253;
assign bias_add_253 = conv_mac_253 + 14'd6579;
logic [31:0] bias_add_254;
assign bias_add_254 = conv_mac_254 + 16'd26550;
logic [31:0] bias_add_255;
assign bias_add_255 = conv_mac_255 + 16'd29925;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[21:15]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[21:15]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[21:15]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[21:15]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[21:15]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[21:15]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[21:15]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[21:15]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[21:15]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[21:15]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[21:15]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[21:15]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[21:15]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[21:15]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[21:15]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[21:15]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[21:15]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[21:15]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[21:15]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[21:15]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[21:15]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[21:15]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[21:15]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[21:15]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[21:15]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[21:15]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[21:15]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[21:15]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[21:15]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[21:15]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[21:15]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[21:15]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[21:15]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[21:15]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[21:15]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[21:15]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[21:15]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[21:15]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[21:15]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[21:15]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[21:15]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[21:15]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[21:15]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[21:15]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[21:15]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[21:15]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[21:15]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[21:15]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[21:15]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[21:15]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[21:15]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[21:15]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[21:15]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[21:15]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[21:15]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[21:15]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[21:15]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[21:15]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[21:15]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[21:15]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[21:15]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[21:15]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[21:15]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[21:15]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[21:15]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[21:15]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[21:15]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[21:15]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[21:15]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[21:15]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[21:15]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[21:15]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[21:15]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[21:15]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[21:15]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[21:15]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[21:15]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[21:15]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[21:15]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[21:15]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[21:15]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[21:15]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[21:15]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[21:15]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[21:15]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[21:15]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[21:15]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[21:15]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[21:15]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[21:15]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[21:15]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[21:15]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[21:15]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[21:15]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[21:15]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[21:15]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[21:15]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[21:15]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[21:15]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[21:15]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[21:15]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[21:15]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[21:15]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[21:15]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[21:15]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[21:15]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[21:15]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[21:15]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[21:15]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[21:15]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[21:15]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[21:15]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[21:15]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[21:15]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[21:15]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[21:15]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[21:15]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[21:15]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[21:15]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[21:15]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[21:15]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[21:15]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[21:15]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[21:15]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[21:15]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[21:15]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[21:15]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[21:15]}} :'d6) : '0;
logic [7:0] relu_128;
assign relu_128[7:0] = (bias_add_128[31]==0) ? ((bias_add_128<3'd6) ? {{bias_add_128[31],bias_add_128[21:15]}} :'d6) : '0;
logic [7:0] relu_129;
assign relu_129[7:0] = (bias_add_129[31]==0) ? ((bias_add_129<3'd6) ? {{bias_add_129[31],bias_add_129[21:15]}} :'d6) : '0;
logic [7:0] relu_130;
assign relu_130[7:0] = (bias_add_130[31]==0) ? ((bias_add_130<3'd6) ? {{bias_add_130[31],bias_add_130[21:15]}} :'d6) : '0;
logic [7:0] relu_131;
assign relu_131[7:0] = (bias_add_131[31]==0) ? ((bias_add_131<3'd6) ? {{bias_add_131[31],bias_add_131[21:15]}} :'d6) : '0;
logic [7:0] relu_132;
assign relu_132[7:0] = (bias_add_132[31]==0) ? ((bias_add_132<3'd6) ? {{bias_add_132[31],bias_add_132[21:15]}} :'d6) : '0;
logic [7:0] relu_133;
assign relu_133[7:0] = (bias_add_133[31]==0) ? ((bias_add_133<3'd6) ? {{bias_add_133[31],bias_add_133[21:15]}} :'d6) : '0;
logic [7:0] relu_134;
assign relu_134[7:0] = (bias_add_134[31]==0) ? ((bias_add_134<3'd6) ? {{bias_add_134[31],bias_add_134[21:15]}} :'d6) : '0;
logic [7:0] relu_135;
assign relu_135[7:0] = (bias_add_135[31]==0) ? ((bias_add_135<3'd6) ? {{bias_add_135[31],bias_add_135[21:15]}} :'d6) : '0;
logic [7:0] relu_136;
assign relu_136[7:0] = (bias_add_136[31]==0) ? ((bias_add_136<3'd6) ? {{bias_add_136[31],bias_add_136[21:15]}} :'d6) : '0;
logic [7:0] relu_137;
assign relu_137[7:0] = (bias_add_137[31]==0) ? ((bias_add_137<3'd6) ? {{bias_add_137[31],bias_add_137[21:15]}} :'d6) : '0;
logic [7:0] relu_138;
assign relu_138[7:0] = (bias_add_138[31]==0) ? ((bias_add_138<3'd6) ? {{bias_add_138[31],bias_add_138[21:15]}} :'d6) : '0;
logic [7:0] relu_139;
assign relu_139[7:0] = (bias_add_139[31]==0) ? ((bias_add_139<3'd6) ? {{bias_add_139[31],bias_add_139[21:15]}} :'d6) : '0;
logic [7:0] relu_140;
assign relu_140[7:0] = (bias_add_140[31]==0) ? ((bias_add_140<3'd6) ? {{bias_add_140[31],bias_add_140[21:15]}} :'d6) : '0;
logic [7:0] relu_141;
assign relu_141[7:0] = (bias_add_141[31]==0) ? ((bias_add_141<3'd6) ? {{bias_add_141[31],bias_add_141[21:15]}} :'d6) : '0;
logic [7:0] relu_142;
assign relu_142[7:0] = (bias_add_142[31]==0) ? ((bias_add_142<3'd6) ? {{bias_add_142[31],bias_add_142[21:15]}} :'d6) : '0;
logic [7:0] relu_143;
assign relu_143[7:0] = (bias_add_143[31]==0) ? ((bias_add_143<3'd6) ? {{bias_add_143[31],bias_add_143[21:15]}} :'d6) : '0;
logic [7:0] relu_144;
assign relu_144[7:0] = (bias_add_144[31]==0) ? ((bias_add_144<3'd6) ? {{bias_add_144[31],bias_add_144[21:15]}} :'d6) : '0;
logic [7:0] relu_145;
assign relu_145[7:0] = (bias_add_145[31]==0) ? ((bias_add_145<3'd6) ? {{bias_add_145[31],bias_add_145[21:15]}} :'d6) : '0;
logic [7:0] relu_146;
assign relu_146[7:0] = (bias_add_146[31]==0) ? ((bias_add_146<3'd6) ? {{bias_add_146[31],bias_add_146[21:15]}} :'d6) : '0;
logic [7:0] relu_147;
assign relu_147[7:0] = (bias_add_147[31]==0) ? ((bias_add_147<3'd6) ? {{bias_add_147[31],bias_add_147[21:15]}} :'d6) : '0;
logic [7:0] relu_148;
assign relu_148[7:0] = (bias_add_148[31]==0) ? ((bias_add_148<3'd6) ? {{bias_add_148[31],bias_add_148[21:15]}} :'d6) : '0;
logic [7:0] relu_149;
assign relu_149[7:0] = (bias_add_149[31]==0) ? ((bias_add_149<3'd6) ? {{bias_add_149[31],bias_add_149[21:15]}} :'d6) : '0;
logic [7:0] relu_150;
assign relu_150[7:0] = (bias_add_150[31]==0) ? ((bias_add_150<3'd6) ? {{bias_add_150[31],bias_add_150[21:15]}} :'d6) : '0;
logic [7:0] relu_151;
assign relu_151[7:0] = (bias_add_151[31]==0) ? ((bias_add_151<3'd6) ? {{bias_add_151[31],bias_add_151[21:15]}} :'d6) : '0;
logic [7:0] relu_152;
assign relu_152[7:0] = (bias_add_152[31]==0) ? ((bias_add_152<3'd6) ? {{bias_add_152[31],bias_add_152[21:15]}} :'d6) : '0;
logic [7:0] relu_153;
assign relu_153[7:0] = (bias_add_153[31]==0) ? ((bias_add_153<3'd6) ? {{bias_add_153[31],bias_add_153[21:15]}} :'d6) : '0;
logic [7:0] relu_154;
assign relu_154[7:0] = (bias_add_154[31]==0) ? ((bias_add_154<3'd6) ? {{bias_add_154[31],bias_add_154[21:15]}} :'d6) : '0;
logic [7:0] relu_155;
assign relu_155[7:0] = (bias_add_155[31]==0) ? ((bias_add_155<3'd6) ? {{bias_add_155[31],bias_add_155[21:15]}} :'d6) : '0;
logic [7:0] relu_156;
assign relu_156[7:0] = (bias_add_156[31]==0) ? ((bias_add_156<3'd6) ? {{bias_add_156[31],bias_add_156[21:15]}} :'d6) : '0;
logic [7:0] relu_157;
assign relu_157[7:0] = (bias_add_157[31]==0) ? ((bias_add_157<3'd6) ? {{bias_add_157[31],bias_add_157[21:15]}} :'d6) : '0;
logic [7:0] relu_158;
assign relu_158[7:0] = (bias_add_158[31]==0) ? ((bias_add_158<3'd6) ? {{bias_add_158[31],bias_add_158[21:15]}} :'d6) : '0;
logic [7:0] relu_159;
assign relu_159[7:0] = (bias_add_159[31]==0) ? ((bias_add_159<3'd6) ? {{bias_add_159[31],bias_add_159[21:15]}} :'d6) : '0;
logic [7:0] relu_160;
assign relu_160[7:0] = (bias_add_160[31]==0) ? ((bias_add_160<3'd6) ? {{bias_add_160[31],bias_add_160[21:15]}} :'d6) : '0;
logic [7:0] relu_161;
assign relu_161[7:0] = (bias_add_161[31]==0) ? ((bias_add_161<3'd6) ? {{bias_add_161[31],bias_add_161[21:15]}} :'d6) : '0;
logic [7:0] relu_162;
assign relu_162[7:0] = (bias_add_162[31]==0) ? ((bias_add_162<3'd6) ? {{bias_add_162[31],bias_add_162[21:15]}} :'d6) : '0;
logic [7:0] relu_163;
assign relu_163[7:0] = (bias_add_163[31]==0) ? ((bias_add_163<3'd6) ? {{bias_add_163[31],bias_add_163[21:15]}} :'d6) : '0;
logic [7:0] relu_164;
assign relu_164[7:0] = (bias_add_164[31]==0) ? ((bias_add_164<3'd6) ? {{bias_add_164[31],bias_add_164[21:15]}} :'d6) : '0;
logic [7:0] relu_165;
assign relu_165[7:0] = (bias_add_165[31]==0) ? ((bias_add_165<3'd6) ? {{bias_add_165[31],bias_add_165[21:15]}} :'d6) : '0;
logic [7:0] relu_166;
assign relu_166[7:0] = (bias_add_166[31]==0) ? ((bias_add_166<3'd6) ? {{bias_add_166[31],bias_add_166[21:15]}} :'d6) : '0;
logic [7:0] relu_167;
assign relu_167[7:0] = (bias_add_167[31]==0) ? ((bias_add_167<3'd6) ? {{bias_add_167[31],bias_add_167[21:15]}} :'d6) : '0;
logic [7:0] relu_168;
assign relu_168[7:0] = (bias_add_168[31]==0) ? ((bias_add_168<3'd6) ? {{bias_add_168[31],bias_add_168[21:15]}} :'d6) : '0;
logic [7:0] relu_169;
assign relu_169[7:0] = (bias_add_169[31]==0) ? ((bias_add_169<3'd6) ? {{bias_add_169[31],bias_add_169[21:15]}} :'d6) : '0;
logic [7:0] relu_170;
assign relu_170[7:0] = (bias_add_170[31]==0) ? ((bias_add_170<3'd6) ? {{bias_add_170[31],bias_add_170[21:15]}} :'d6) : '0;
logic [7:0] relu_171;
assign relu_171[7:0] = (bias_add_171[31]==0) ? ((bias_add_171<3'd6) ? {{bias_add_171[31],bias_add_171[21:15]}} :'d6) : '0;
logic [7:0] relu_172;
assign relu_172[7:0] = (bias_add_172[31]==0) ? ((bias_add_172<3'd6) ? {{bias_add_172[31],bias_add_172[21:15]}} :'d6) : '0;
logic [7:0] relu_173;
assign relu_173[7:0] = (bias_add_173[31]==0) ? ((bias_add_173<3'd6) ? {{bias_add_173[31],bias_add_173[21:15]}} :'d6) : '0;
logic [7:0] relu_174;
assign relu_174[7:0] = (bias_add_174[31]==0) ? ((bias_add_174<3'd6) ? {{bias_add_174[31],bias_add_174[21:15]}} :'d6) : '0;
logic [7:0] relu_175;
assign relu_175[7:0] = (bias_add_175[31]==0) ? ((bias_add_175<3'd6) ? {{bias_add_175[31],bias_add_175[21:15]}} :'d6) : '0;
logic [7:0] relu_176;
assign relu_176[7:0] = (bias_add_176[31]==0) ? ((bias_add_176<3'd6) ? {{bias_add_176[31],bias_add_176[21:15]}} :'d6) : '0;
logic [7:0] relu_177;
assign relu_177[7:0] = (bias_add_177[31]==0) ? ((bias_add_177<3'd6) ? {{bias_add_177[31],bias_add_177[21:15]}} :'d6) : '0;
logic [7:0] relu_178;
assign relu_178[7:0] = (bias_add_178[31]==0) ? ((bias_add_178<3'd6) ? {{bias_add_178[31],bias_add_178[21:15]}} :'d6) : '0;
logic [7:0] relu_179;
assign relu_179[7:0] = (bias_add_179[31]==0) ? ((bias_add_179<3'd6) ? {{bias_add_179[31],bias_add_179[21:15]}} :'d6) : '0;
logic [7:0] relu_180;
assign relu_180[7:0] = (bias_add_180[31]==0) ? ((bias_add_180<3'd6) ? {{bias_add_180[31],bias_add_180[21:15]}} :'d6) : '0;
logic [7:0] relu_181;
assign relu_181[7:0] = (bias_add_181[31]==0) ? ((bias_add_181<3'd6) ? {{bias_add_181[31],bias_add_181[21:15]}} :'d6) : '0;
logic [7:0] relu_182;
assign relu_182[7:0] = (bias_add_182[31]==0) ? ((bias_add_182<3'd6) ? {{bias_add_182[31],bias_add_182[21:15]}} :'d6) : '0;
logic [7:0] relu_183;
assign relu_183[7:0] = (bias_add_183[31]==0) ? ((bias_add_183<3'd6) ? {{bias_add_183[31],bias_add_183[21:15]}} :'d6) : '0;
logic [7:0] relu_184;
assign relu_184[7:0] = (bias_add_184[31]==0) ? ((bias_add_184<3'd6) ? {{bias_add_184[31],bias_add_184[21:15]}} :'d6) : '0;
logic [7:0] relu_185;
assign relu_185[7:0] = (bias_add_185[31]==0) ? ((bias_add_185<3'd6) ? {{bias_add_185[31],bias_add_185[21:15]}} :'d6) : '0;
logic [7:0] relu_186;
assign relu_186[7:0] = (bias_add_186[31]==0) ? ((bias_add_186<3'd6) ? {{bias_add_186[31],bias_add_186[21:15]}} :'d6) : '0;
logic [7:0] relu_187;
assign relu_187[7:0] = (bias_add_187[31]==0) ? ((bias_add_187<3'd6) ? {{bias_add_187[31],bias_add_187[21:15]}} :'d6) : '0;
logic [7:0] relu_188;
assign relu_188[7:0] = (bias_add_188[31]==0) ? ((bias_add_188<3'd6) ? {{bias_add_188[31],bias_add_188[21:15]}} :'d6) : '0;
logic [7:0] relu_189;
assign relu_189[7:0] = (bias_add_189[31]==0) ? ((bias_add_189<3'd6) ? {{bias_add_189[31],bias_add_189[21:15]}} :'d6) : '0;
logic [7:0] relu_190;
assign relu_190[7:0] = (bias_add_190[31]==0) ? ((bias_add_190<3'd6) ? {{bias_add_190[31],bias_add_190[21:15]}} :'d6) : '0;
logic [7:0] relu_191;
assign relu_191[7:0] = (bias_add_191[31]==0) ? ((bias_add_191<3'd6) ? {{bias_add_191[31],bias_add_191[21:15]}} :'d6) : '0;
logic [7:0] relu_192;
assign relu_192[7:0] = (bias_add_192[31]==0) ? ((bias_add_192<3'd6) ? {{bias_add_192[31],bias_add_192[21:15]}} :'d6) : '0;
logic [7:0] relu_193;
assign relu_193[7:0] = (bias_add_193[31]==0) ? ((bias_add_193<3'd6) ? {{bias_add_193[31],bias_add_193[21:15]}} :'d6) : '0;
logic [7:0] relu_194;
assign relu_194[7:0] = (bias_add_194[31]==0) ? ((bias_add_194<3'd6) ? {{bias_add_194[31],bias_add_194[21:15]}} :'d6) : '0;
logic [7:0] relu_195;
assign relu_195[7:0] = (bias_add_195[31]==0) ? ((bias_add_195<3'd6) ? {{bias_add_195[31],bias_add_195[21:15]}} :'d6) : '0;
logic [7:0] relu_196;
assign relu_196[7:0] = (bias_add_196[31]==0) ? ((bias_add_196<3'd6) ? {{bias_add_196[31],bias_add_196[21:15]}} :'d6) : '0;
logic [7:0] relu_197;
assign relu_197[7:0] = (bias_add_197[31]==0) ? ((bias_add_197<3'd6) ? {{bias_add_197[31],bias_add_197[21:15]}} :'d6) : '0;
logic [7:0] relu_198;
assign relu_198[7:0] = (bias_add_198[31]==0) ? ((bias_add_198<3'd6) ? {{bias_add_198[31],bias_add_198[21:15]}} :'d6) : '0;
logic [7:0] relu_199;
assign relu_199[7:0] = (bias_add_199[31]==0) ? ((bias_add_199<3'd6) ? {{bias_add_199[31],bias_add_199[21:15]}} :'d6) : '0;
logic [7:0] relu_200;
assign relu_200[7:0] = (bias_add_200[31]==0) ? ((bias_add_200<3'd6) ? {{bias_add_200[31],bias_add_200[21:15]}} :'d6) : '0;
logic [7:0] relu_201;
assign relu_201[7:0] = (bias_add_201[31]==0) ? ((bias_add_201<3'd6) ? {{bias_add_201[31],bias_add_201[21:15]}} :'d6) : '0;
logic [7:0] relu_202;
assign relu_202[7:0] = (bias_add_202[31]==0) ? ((bias_add_202<3'd6) ? {{bias_add_202[31],bias_add_202[21:15]}} :'d6) : '0;
logic [7:0] relu_203;
assign relu_203[7:0] = (bias_add_203[31]==0) ? ((bias_add_203<3'd6) ? {{bias_add_203[31],bias_add_203[21:15]}} :'d6) : '0;
logic [7:0] relu_204;
assign relu_204[7:0] = (bias_add_204[31]==0) ? ((bias_add_204<3'd6) ? {{bias_add_204[31],bias_add_204[21:15]}} :'d6) : '0;
logic [7:0] relu_205;
assign relu_205[7:0] = (bias_add_205[31]==0) ? ((bias_add_205<3'd6) ? {{bias_add_205[31],bias_add_205[21:15]}} :'d6) : '0;
logic [7:0] relu_206;
assign relu_206[7:0] = (bias_add_206[31]==0) ? ((bias_add_206<3'd6) ? {{bias_add_206[31],bias_add_206[21:15]}} :'d6) : '0;
logic [7:0] relu_207;
assign relu_207[7:0] = (bias_add_207[31]==0) ? ((bias_add_207<3'd6) ? {{bias_add_207[31],bias_add_207[21:15]}} :'d6) : '0;
logic [7:0] relu_208;
assign relu_208[7:0] = (bias_add_208[31]==0) ? ((bias_add_208<3'd6) ? {{bias_add_208[31],bias_add_208[21:15]}} :'d6) : '0;
logic [7:0] relu_209;
assign relu_209[7:0] = (bias_add_209[31]==0) ? ((bias_add_209<3'd6) ? {{bias_add_209[31],bias_add_209[21:15]}} :'d6) : '0;
logic [7:0] relu_210;
assign relu_210[7:0] = (bias_add_210[31]==0) ? ((bias_add_210<3'd6) ? {{bias_add_210[31],bias_add_210[21:15]}} :'d6) : '0;
logic [7:0] relu_211;
assign relu_211[7:0] = (bias_add_211[31]==0) ? ((bias_add_211<3'd6) ? {{bias_add_211[31],bias_add_211[21:15]}} :'d6) : '0;
logic [7:0] relu_212;
assign relu_212[7:0] = (bias_add_212[31]==0) ? ((bias_add_212<3'd6) ? {{bias_add_212[31],bias_add_212[21:15]}} :'d6) : '0;
logic [7:0] relu_213;
assign relu_213[7:0] = (bias_add_213[31]==0) ? ((bias_add_213<3'd6) ? {{bias_add_213[31],bias_add_213[21:15]}} :'d6) : '0;
logic [7:0] relu_214;
assign relu_214[7:0] = (bias_add_214[31]==0) ? ((bias_add_214<3'd6) ? {{bias_add_214[31],bias_add_214[21:15]}} :'d6) : '0;
logic [7:0] relu_215;
assign relu_215[7:0] = (bias_add_215[31]==0) ? ((bias_add_215<3'd6) ? {{bias_add_215[31],bias_add_215[21:15]}} :'d6) : '0;
logic [7:0] relu_216;
assign relu_216[7:0] = (bias_add_216[31]==0) ? ((bias_add_216<3'd6) ? {{bias_add_216[31],bias_add_216[21:15]}} :'d6) : '0;
logic [7:0] relu_217;
assign relu_217[7:0] = (bias_add_217[31]==0) ? ((bias_add_217<3'd6) ? {{bias_add_217[31],bias_add_217[21:15]}} :'d6) : '0;
logic [7:0] relu_218;
assign relu_218[7:0] = (bias_add_218[31]==0) ? ((bias_add_218<3'd6) ? {{bias_add_218[31],bias_add_218[21:15]}} :'d6) : '0;
logic [7:0] relu_219;
assign relu_219[7:0] = (bias_add_219[31]==0) ? ((bias_add_219<3'd6) ? {{bias_add_219[31],bias_add_219[21:15]}} :'d6) : '0;
logic [7:0] relu_220;
assign relu_220[7:0] = (bias_add_220[31]==0) ? ((bias_add_220<3'd6) ? {{bias_add_220[31],bias_add_220[21:15]}} :'d6) : '0;
logic [7:0] relu_221;
assign relu_221[7:0] = (bias_add_221[31]==0) ? ((bias_add_221<3'd6) ? {{bias_add_221[31],bias_add_221[21:15]}} :'d6) : '0;
logic [7:0] relu_222;
assign relu_222[7:0] = (bias_add_222[31]==0) ? ((bias_add_222<3'd6) ? {{bias_add_222[31],bias_add_222[21:15]}} :'d6) : '0;
logic [7:0] relu_223;
assign relu_223[7:0] = (bias_add_223[31]==0) ? ((bias_add_223<3'd6) ? {{bias_add_223[31],bias_add_223[21:15]}} :'d6) : '0;
logic [7:0] relu_224;
assign relu_224[7:0] = (bias_add_224[31]==0) ? ((bias_add_224<3'd6) ? {{bias_add_224[31],bias_add_224[21:15]}} :'d6) : '0;
logic [7:0] relu_225;
assign relu_225[7:0] = (bias_add_225[31]==0) ? ((bias_add_225<3'd6) ? {{bias_add_225[31],bias_add_225[21:15]}} :'d6) : '0;
logic [7:0] relu_226;
assign relu_226[7:0] = (bias_add_226[31]==0) ? ((bias_add_226<3'd6) ? {{bias_add_226[31],bias_add_226[21:15]}} :'d6) : '0;
logic [7:0] relu_227;
assign relu_227[7:0] = (bias_add_227[31]==0) ? ((bias_add_227<3'd6) ? {{bias_add_227[31],bias_add_227[21:15]}} :'d6) : '0;
logic [7:0] relu_228;
assign relu_228[7:0] = (bias_add_228[31]==0) ? ((bias_add_228<3'd6) ? {{bias_add_228[31],bias_add_228[21:15]}} :'d6) : '0;
logic [7:0] relu_229;
assign relu_229[7:0] = (bias_add_229[31]==0) ? ((bias_add_229<3'd6) ? {{bias_add_229[31],bias_add_229[21:15]}} :'d6) : '0;
logic [7:0] relu_230;
assign relu_230[7:0] = (bias_add_230[31]==0) ? ((bias_add_230<3'd6) ? {{bias_add_230[31],bias_add_230[21:15]}} :'d6) : '0;
logic [7:0] relu_231;
assign relu_231[7:0] = (bias_add_231[31]==0) ? ((bias_add_231<3'd6) ? {{bias_add_231[31],bias_add_231[21:15]}} :'d6) : '0;
logic [7:0] relu_232;
assign relu_232[7:0] = (bias_add_232[31]==0) ? ((bias_add_232<3'd6) ? {{bias_add_232[31],bias_add_232[21:15]}} :'d6) : '0;
logic [7:0] relu_233;
assign relu_233[7:0] = (bias_add_233[31]==0) ? ((bias_add_233<3'd6) ? {{bias_add_233[31],bias_add_233[21:15]}} :'d6) : '0;
logic [7:0] relu_234;
assign relu_234[7:0] = (bias_add_234[31]==0) ? ((bias_add_234<3'd6) ? {{bias_add_234[31],bias_add_234[21:15]}} :'d6) : '0;
logic [7:0] relu_235;
assign relu_235[7:0] = (bias_add_235[31]==0) ? ((bias_add_235<3'd6) ? {{bias_add_235[31],bias_add_235[21:15]}} :'d6) : '0;
logic [7:0] relu_236;
assign relu_236[7:0] = (bias_add_236[31]==0) ? ((bias_add_236<3'd6) ? {{bias_add_236[31],bias_add_236[21:15]}} :'d6) : '0;
logic [7:0] relu_237;
assign relu_237[7:0] = (bias_add_237[31]==0) ? ((bias_add_237<3'd6) ? {{bias_add_237[31],bias_add_237[21:15]}} :'d6) : '0;
logic [7:0] relu_238;
assign relu_238[7:0] = (bias_add_238[31]==0) ? ((bias_add_238<3'd6) ? {{bias_add_238[31],bias_add_238[21:15]}} :'d6) : '0;
logic [7:0] relu_239;
assign relu_239[7:0] = (bias_add_239[31]==0) ? ((bias_add_239<3'd6) ? {{bias_add_239[31],bias_add_239[21:15]}} :'d6) : '0;
logic [7:0] relu_240;
assign relu_240[7:0] = (bias_add_240[31]==0) ? ((bias_add_240<3'd6) ? {{bias_add_240[31],bias_add_240[21:15]}} :'d6) : '0;
logic [7:0] relu_241;
assign relu_241[7:0] = (bias_add_241[31]==0) ? ((bias_add_241<3'd6) ? {{bias_add_241[31],bias_add_241[21:15]}} :'d6) : '0;
logic [7:0] relu_242;
assign relu_242[7:0] = (bias_add_242[31]==0) ? ((bias_add_242<3'd6) ? {{bias_add_242[31],bias_add_242[21:15]}} :'d6) : '0;
logic [7:0] relu_243;
assign relu_243[7:0] = (bias_add_243[31]==0) ? ((bias_add_243<3'd6) ? {{bias_add_243[31],bias_add_243[21:15]}} :'d6) : '0;
logic [7:0] relu_244;
assign relu_244[7:0] = (bias_add_244[31]==0) ? ((bias_add_244<3'd6) ? {{bias_add_244[31],bias_add_244[21:15]}} :'d6) : '0;
logic [7:0] relu_245;
assign relu_245[7:0] = (bias_add_245[31]==0) ? ((bias_add_245<3'd6) ? {{bias_add_245[31],bias_add_245[21:15]}} :'d6) : '0;
logic [7:0] relu_246;
assign relu_246[7:0] = (bias_add_246[31]==0) ? ((bias_add_246<3'd6) ? {{bias_add_246[31],bias_add_246[21:15]}} :'d6) : '0;
logic [7:0] relu_247;
assign relu_247[7:0] = (bias_add_247[31]==0) ? ((bias_add_247<3'd6) ? {{bias_add_247[31],bias_add_247[21:15]}} :'d6) : '0;
logic [7:0] relu_248;
assign relu_248[7:0] = (bias_add_248[31]==0) ? ((bias_add_248<3'd6) ? {{bias_add_248[31],bias_add_248[21:15]}} :'d6) : '0;
logic [7:0] relu_249;
assign relu_249[7:0] = (bias_add_249[31]==0) ? ((bias_add_249<3'd6) ? {{bias_add_249[31],bias_add_249[21:15]}} :'d6) : '0;
logic [7:0] relu_250;
assign relu_250[7:0] = (bias_add_250[31]==0) ? ((bias_add_250<3'd6) ? {{bias_add_250[31],bias_add_250[21:15]}} :'d6) : '0;
logic [7:0] relu_251;
assign relu_251[7:0] = (bias_add_251[31]==0) ? ((bias_add_251<3'd6) ? {{bias_add_251[31],bias_add_251[21:15]}} :'d6) : '0;
logic [7:0] relu_252;
assign relu_252[7:0] = (bias_add_252[31]==0) ? ((bias_add_252<3'd6) ? {{bias_add_252[31],bias_add_252[21:15]}} :'d6) : '0;
logic [7:0] relu_253;
assign relu_253[7:0] = (bias_add_253[31]==0) ? ((bias_add_253<3'd6) ? {{bias_add_253[31],bias_add_253[21:15]}} :'d6) : '0;
logic [7:0] relu_254;
assign relu_254[7:0] = (bias_add_254[31]==0) ? ((bias_add_254<3'd6) ? {{bias_add_254[31],bias_add_254[21:15]}} :'d6) : '0;
logic [7:0] relu_255;
assign relu_255[7:0] = (bias_add_255[31]==0) ? ((bias_add_255<3'd6) ? {{bias_add_255[31],bias_add_255[21:15]}} :'d6) : '0;

assign output_act = {
	relu_255,
	relu_254,
	relu_253,
	relu_252,
	relu_251,
	relu_250,
	relu_249,
	relu_248,
	relu_247,
	relu_246,
	relu_245,
	relu_244,
	relu_243,
	relu_242,
	relu_241,
	relu_240,
	relu_239,
	relu_238,
	relu_237,
	relu_236,
	relu_235,
	relu_234,
	relu_233,
	relu_232,
	relu_231,
	relu_230,
	relu_229,
	relu_228,
	relu_227,
	relu_226,
	relu_225,
	relu_224,
	relu_223,
	relu_222,
	relu_221,
	relu_220,
	relu_219,
	relu_218,
	relu_217,
	relu_216,
	relu_215,
	relu_214,
	relu_213,
	relu_212,
	relu_211,
	relu_210,
	relu_209,
	relu_208,
	relu_207,
	relu_206,
	relu_205,
	relu_204,
	relu_203,
	relu_202,
	relu_201,
	relu_200,
	relu_199,
	relu_198,
	relu_197,
	relu_196,
	relu_195,
	relu_194,
	relu_193,
	relu_192,
	relu_191,
	relu_190,
	relu_189,
	relu_188,
	relu_187,
	relu_186,
	relu_185,
	relu_184,
	relu_183,
	relu_182,
	relu_181,
	relu_180,
	relu_179,
	relu_178,
	relu_177,
	relu_176,
	relu_175,
	relu_174,
	relu_173,
	relu_172,
	relu_171,
	relu_170,
	relu_169,
	relu_168,
	relu_167,
	relu_166,
	relu_165,
	relu_164,
	relu_163,
	relu_162,
	relu_161,
	relu_160,
	relu_159,
	relu_158,
	relu_157,
	relu_156,
	relu_155,
	relu_154,
	relu_153,
	relu_152,
	relu_151,
	relu_150,
	relu_149,
	relu_148,
	relu_147,
	relu_146,
	relu_145,
	relu_144,
	relu_143,
	relu_142,
	relu_141,
	relu_140,
	relu_139,
	relu_138,
	relu_137,
	relu_136,
	relu_135,
	relu_134,
	relu_133,
	relu_132,
	relu_131,
	relu_130,
	relu_129,
	relu_128,
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
