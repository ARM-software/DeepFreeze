module conv11_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [1024-1:0] input_act,
    output logic [1024-1:0] output_act,
    output logic ready
);

logic [1024-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 15'sd 10068) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20766) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1729) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_6[7:0]) +
	( 11'sd 806) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6760) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7896) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15748) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16007) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18534) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25282) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25733) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1090) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25385) * $signed(input_fmap_23[7:0]) +
	( 11'sd 774) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1152) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20236) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6078) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16931) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6847) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20090) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30974) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1671) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10473) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13461) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23303) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18755) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2657) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32499) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1806) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12495) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29242) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19871) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29758) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2090) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3383) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16271) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14670) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13638) * $signed(input_fmap_61[7:0]) +
	( 8'sd 109) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27842) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29151) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21737) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15647) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3737) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14903) * $signed(input_fmap_72[7:0]) +
	( 10'sd 477) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23046) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8787) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2176) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22090) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21706) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15982) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11405) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16999) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16432) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29505) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_88[7:0]) +
	( 10'sd 500) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20604) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30904) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32072) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_96[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15939) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2267) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16213) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19112) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8243) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12212) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32648) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22727) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19810) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10819) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19662) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13979) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1075) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11761) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30652) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 15'sd 10209) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25495) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6300) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27449) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14371) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17099) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29126) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29013) * $signed(input_fmap_9[7:0]) +
	( 13'sd 4079) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10041) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10086) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19462) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30862) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19596) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12289) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7368) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6107) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11594) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5778) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19705) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12378) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25858) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_33[7:0]) +
	( 10'sd 490) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10902) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14489) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9791) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23783) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24605) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9614) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13652) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17189) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11230) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19214) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32365) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29469) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29878) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19812) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30157) * $signed(input_fmap_57[7:0]) +
	( 9'sd 245) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17229) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13855) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12116) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8622) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4998) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8262) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25840) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24057) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13442) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10532) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11842) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28663) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30299) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1209) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12030) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31529) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4844) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14403) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_86[7:0]) +
	( 11'sd 768) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16449) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25065) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17666) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9608) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11418) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19782) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14587) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13738) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30082) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2671) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20866) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2720) * $signed(input_fmap_106[7:0]) +
	( 10'sd 447) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5864) * $signed(input_fmap_108[7:0]) +
	( 11'sd 1002) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20114) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26266) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6013) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9299) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11660) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9530) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25016) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16408) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3712) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26217) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 15'sd 13275) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15525) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7427) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23617) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23671) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21287) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14205) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20321) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4840) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10387) * $signed(input_fmap_16[7:0]) +
	( 10'sd 334) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8629) * $signed(input_fmap_18[7:0]) +
	( 11'sd 589) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28760) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14206) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2814) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26615) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15759) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13864) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5001) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28517) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10149) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21225) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16326) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31537) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18170) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9648) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28408) * $signed(input_fmap_40[7:0]) +
	( 11'sd 642) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20227) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28270) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4392) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1641) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18813) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32217) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16384) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17278) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29895) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3555) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30572) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8234) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20079) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10707) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20832) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10917) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21208) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1234) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21228) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22475) * $signed(input_fmap_76[7:0]) +
	( 11'sd 899) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24768) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28413) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30706) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17337) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17276) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10784) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20442) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7761) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15863) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29448) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11823) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14548) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10637) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9546) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4361) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2942) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19426) * $signed(input_fmap_104[7:0]) +
	( 11'sd 673) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20714) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30190) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21798) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3630) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6217) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27910) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31225) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10790) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8470) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17153) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1086) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26173) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14340) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29540) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 14'sd 5603) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6159) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27776) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1652) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9357) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20170) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15205) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12538) * $signed(input_fmap_11[7:0]) +
	( 7'sd 51) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23741) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16803) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26772) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31291) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20538) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21025) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9654) * $signed(input_fmap_24[7:0]) +
	( 10'sd 268) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29899) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25691) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27620) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1114) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17398) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17226) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24584) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19022) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26231) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6727) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14916) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18589) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32363) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24378) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12131) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20785) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9707) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20934) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28006) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19352) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8663) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14082) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12707) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27254) * $signed(input_fmap_62[7:0]) +
	( 11'sd 548) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27300) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11100) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11648) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11410) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_71[7:0]) +
	( 13'sd 4049) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2566) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8994) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11066) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2096) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20597) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25780) * $signed(input_fmap_83[7:0]) +
	( 11'sd 798) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18847) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6897) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6954) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20461) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30891) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19134) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23904) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29943) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17915) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25896) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22391) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29443) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17756) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24115) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13061) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3294) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27731) * $signed(input_fmap_109[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31840) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10980) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2692) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3397) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19208) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10022) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6320) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21083) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24040) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31497) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4667) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9234) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24750) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1675) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 16'sd 18675) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17363) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12970) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16531) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12887) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7227) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23298) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28444) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24633) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21228) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7300) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26337) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24462) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3602) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12704) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3976) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2367) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18740) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6633) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28065) * $signed(input_fmap_20[7:0]) +
	( 11'sd 715) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30662) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11590) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2209) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22320) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3286) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29054) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12538) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31972) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30881) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16604) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16076) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17093) * $signed(input_fmap_42[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13319) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7617) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2053) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20626) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27849) * $signed(input_fmap_55[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9378) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1216) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25229) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17623) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21631) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25360) * $signed(input_fmap_71[7:0]) +
	( 9'sd 253) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22256) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2624) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10198) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28006) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8419) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5293) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28512) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27074) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10273) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9305) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13555) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18690) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3448) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30129) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30393) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5250) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_100[7:0]) +
	( 10'sd 412) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12397) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31410) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4128) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13575) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27422) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10086) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15876) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11748) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18401) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8552) * $signed(input_fmap_114[7:0]) +
	( 11'sd 529) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32303) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8088) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17959) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23454) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18552) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29326) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7538) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20518) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10364) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 16'sd 31552) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5760) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5096) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27883) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12298) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21855) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26431) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19411) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23780) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11945) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32383) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19088) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25077) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31864) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26012) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9144) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4817) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32522) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19482) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23272) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32633) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4763) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6522) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13869) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30611) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9004) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31733) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1331) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26628) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20118) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1580) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31134) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4342) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23311) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1884) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6600) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26334) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14926) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14404) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7784) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32368) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13446) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21400) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29862) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17892) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5023) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14517) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23207) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28847) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10587) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12830) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26448) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3021) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19674) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18904) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25534) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16637) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3678) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5054) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7805) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24504) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13708) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13818) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7795) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7086) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26661) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28476) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12189) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2734) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13631) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6730) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11409) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17741) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30047) * $signed(input_fmap_114[7:0]) +
	( 10'sd 389) * $signed(input_fmap_115[7:0]) +
	( 11'sd 808) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20588) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25434) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8590) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18420) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6980) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31701) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19523) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20331) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 15'sd 9354) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12438) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1345) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8838) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17240) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7476) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11112) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2055) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27312) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6915) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_16[7:0]) +
	( 11'sd 879) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23749) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2389) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9385) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13926) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6080) * $signed(input_fmap_24[7:0]) +
	( 13'sd 4008) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32473) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12065) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29425) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24931) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23789) * $signed(input_fmap_30[7:0]) +
	( 11'sd 800) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21523) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32201) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29805) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7824) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32589) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12785) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27329) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16636) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8366) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_54[7:0]) +
	( 11'sd 711) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2523) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13488) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24495) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14068) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5435) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23822) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_64[7:0]) +
	( 11'sd 858) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2449) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23290) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13095) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11750) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25858) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7061) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9188) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4534) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26397) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8060) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11100) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25314) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23788) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1407) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11202) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25920) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16080) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9949) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6223) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21760) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32037) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26019) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15216) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18107) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16707) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8585) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_104[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12153) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18278) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30925) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16123) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15444) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4482) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_113[7:0]) +
	( 6'sd 20) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_115[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26611) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29210) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1516) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27913) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4742) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29208) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31245) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11313) * $signed(input_fmap_125[7:0]) +
	( 11'sd 682) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14449) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 11'sd 610) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29453) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7851) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15289) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19569) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21292) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20112) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31102) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20118) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23662) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19542) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20954) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13385) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6570) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1603) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2301) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25473) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24125) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15372) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29063) * $signed(input_fmap_26[7:0]) +
	( 10'sd 444) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30846) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31234) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12339) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18834) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15352) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2553) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22159) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16509) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14610) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13693) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14185) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3226) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21357) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1730) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12016) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19023) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28465) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8099) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12580) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7045) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12751) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5085) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18015) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9350) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22275) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11125) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7081) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25501) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27487) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22983) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15904) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19324) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13699) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4123) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_86[7:0]) +
	( 8'sd 75) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4383) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4113) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19624) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13950) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22820) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14447) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1620) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_99[7:0]) +
	( 10'sd 293) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_104[7:0]) +
	( 11'sd 859) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9488) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20853) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2248) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4788) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31127) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3060) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12724) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5341) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24934) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12266) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9968) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28376) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 16'sd 30927) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22372) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15017) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5141) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20115) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19681) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23032) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7528) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26165) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22822) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27019) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13477) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21068) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22486) * $signed(input_fmap_16[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9546) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2184) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15015) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20718) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22426) * $signed(input_fmap_22[7:0]) +
	( 11'sd 600) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20474) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32174) * $signed(input_fmap_26[7:0]) +
	( 11'sd 830) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24764) * $signed(input_fmap_28[7:0]) +
	( 11'sd 995) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16212) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17994) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19020) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17566) * $signed(input_fmap_35[7:0]) +
	( 5'sd 15) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16092) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29914) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21177) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14842) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14451) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5559) * $signed(input_fmap_47[7:0]) +
	( 14'sd 8033) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26813) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21419) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30826) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10943) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30849) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16376) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5452) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1947) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14222) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28106) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28029) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17452) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15572) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23076) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7506) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13388) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20436) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21060) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5580) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16821) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4318) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7762) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12847) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26584) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31632) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14478) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6745) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10968) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17261) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8354) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28234) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10677) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26945) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22707) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17822) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28502) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29755) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9970) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12383) * $signed(input_fmap_106[7:0]) +
	( 10'sd 363) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18680) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32692) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28711) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23944) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25787) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22373) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10608) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31144) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17995) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30352) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26874) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2714) * $signed(input_fmap_125[7:0]) +
	( 11'sd 677) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 16'sd 32454) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20359) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31832) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30583) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3863) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21836) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10839) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4752) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17691) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32273) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15561) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8566) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2129) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12665) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1173) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30387) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17881) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27802) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5308) * $signed(input_fmap_28[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9870) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26551) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6146) * $signed(input_fmap_33[7:0]) +
	( 11'sd 557) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10411) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16932) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7362) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18427) * $signed(input_fmap_43[7:0]) +
	( 11'sd 569) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7618) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24165) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23522) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2366) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26763) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18821) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14474) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15299) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12440) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2306) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11341) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29005) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24076) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31827) * $signed(input_fmap_67[7:0]) +
	( 10'sd 445) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27188) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13351) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32365) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22584) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29220) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32368) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28962) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5436) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14893) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26881) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14573) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20121) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8576) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14006) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6357) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1828) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9280) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10492) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28745) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20124) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2300) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24077) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17150) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6665) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30286) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13207) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23837) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12209) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6125) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6518) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15583) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13567) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19629) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1076) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24646) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15400) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2822) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9440) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26822) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3768) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18671) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 16'sd 31523) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25527) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17931) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21818) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11560) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7148) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20692) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13513) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32396) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26154) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23834) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23272) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2053) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6278) * $signed(input_fmap_23[7:0]) +
	( 11'sd 589) * $signed(input_fmap_24[7:0]) +
	( 11'sd 1000) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7622) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30867) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7950) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4637) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27048) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19080) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17712) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18729) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4523) * $signed(input_fmap_38[7:0]) +
	( 10'sd 297) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24765) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32523) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12916) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16346) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7391) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19942) * $signed(input_fmap_48[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8977) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23208) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_52[7:0]) +
	( 11'sd 996) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24373) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17000) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32136) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32028) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6881) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5402) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31465) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22355) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15553) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32249) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7293) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18082) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21990) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1876) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10860) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15133) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26250) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21140) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24056) * $signed(input_fmap_77[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1497) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18592) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31568) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5947) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4374) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9463) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27047) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22561) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9449) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16783) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9897) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15327) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28081) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21363) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9352) * $signed(input_fmap_102[7:0]) +
	( 10'sd 423) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32060) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21434) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22863) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21862) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5606) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30588) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7473) * $signed(input_fmap_114[7:0]) +
	( 11'sd 587) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2079) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20300) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1507) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_119[7:0]) +
	( 11'sd 854) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11261) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29756) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22153) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8407) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 16'sd 31612) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15723) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8453) * $signed(input_fmap_6[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_8[7:0]) +
	( 13'sd 4071) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1120) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30979) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16699) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_15[7:0]) +
	( 11'sd 910) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15245) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14566) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17716) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25767) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4477) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2643) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20456) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30514) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20535) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22378) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20786) * $signed(input_fmap_33[7:0]) +
	( 9'sd 149) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27387) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3454) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1262) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14430) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29192) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_43[7:0]) +
	( 10'sd 397) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7470) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15381) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29930) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21388) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23948) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3879) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21550) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21583) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24509) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8263) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18708) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11413) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24575) * $signed(input_fmap_63[7:0]) +
	( 11'sd 979) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20859) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5300) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15036) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19124) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20966) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19651) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19361) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24667) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20815) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14557) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1156) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29794) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11732) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15557) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16305) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7899) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16089) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26431) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12690) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32357) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31616) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3031) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28658) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31379) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27351) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1066) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15158) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29880) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27919) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22908) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21737) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15282) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30147) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2515) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16007) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11380) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10018) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1107) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5586) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4521) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 12'sd 1036) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10784) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30501) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29105) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25337) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15608) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10013) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7847) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31396) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28591) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17110) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32558) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8675) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17029) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16331) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21529) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13034) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9703) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13862) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23064) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7573) * $signed(input_fmap_34[7:0]) +
	( 9'sd 138) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21430) * $signed(input_fmap_37[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22450) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19581) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29412) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29996) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10972) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4445) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29820) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15896) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24307) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12594) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4207) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18347) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21097) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1166) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32524) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32716) * $signed(input_fmap_64[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5704) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9085) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26234) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29414) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4940) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6472) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23759) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15003) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9031) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6818) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29956) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26574) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30071) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19351) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10011) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4308) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30162) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7032) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8973) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9559) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30762) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2767) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14558) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31968) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11453) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12253) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26673) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22245) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24736) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13688) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_110[7:0]) +
	( 11'sd 798) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4200) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_115[7:0]) +
	( 11'sd 727) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2777) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8964) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_122[7:0]) +
	( 11'sd 585) * $signed(input_fmap_123[7:0]) +
	( 10'sd 466) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16951) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20720) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 16'sd 17783) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10829) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24032) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29028) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5697) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30957) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30667) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6653) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17494) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21299) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13787) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25427) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5223) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4949) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7801) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28413) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26591) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16400) * $signed(input_fmap_24[7:0]) +
	( 9'sd 139) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9547) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28156) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14773) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16951) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1844) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2753) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7092) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2955) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8255) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26766) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11490) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8310) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29521) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26883) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14289) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17142) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6199) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3841) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23191) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9179) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19230) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25049) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12100) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22704) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18183) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27701) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23866) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5292) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29382) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19251) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14246) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30326) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20381) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24471) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2456) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25806) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16145) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4676) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11146) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13582) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14294) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10663) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32583) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25180) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5536) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15601) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14403) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23083) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24017) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12107) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12846) * $signed(input_fmap_100[7:0]) +
	( 11'sd 655) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27931) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26791) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25971) * $signed(input_fmap_106[7:0]) +
	( 13'sd 4053) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21552) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7425) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22419) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1829) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18652) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28309) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19884) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2791) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7710) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7673) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26461) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_121[7:0]) +
	( 8'sd 119) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23207) * $signed(input_fmap_125[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26810) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 16'sd 17551) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8070) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16393) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22418) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22475) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15537) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12705) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18672) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13594) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16330) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27388) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31330) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14385) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29771) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21738) * $signed(input_fmap_23[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7588) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30371) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24091) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20058) * $signed(input_fmap_30[7:0]) +
	( 11'sd 567) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2573) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15372) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3122) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19548) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21681) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1189) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1891) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22773) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28465) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19056) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2849) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23637) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1914) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9948) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11371) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30360) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23748) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28070) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9736) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5662) * $signed(input_fmap_59[7:0]) +
	( 9'sd 198) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3936) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22640) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12233) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26542) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16340) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6747) * $signed(input_fmap_68[7:0]) +
	( 9'sd 228) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2744) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28857) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23814) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13901) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2405) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15844) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13777) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21181) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9858) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11675) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8974) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1951) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17738) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5985) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22766) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17693) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12032) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28978) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19252) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1221) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23752) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29411) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2436) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11702) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12301) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4726) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32198) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13257) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8552) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8598) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24178) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22292) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30460) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10687) * $signed(input_fmap_123[7:0]) +
	( 11'sd 630) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10425) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13913) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 14'sd 6578) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21529) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15394) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14220) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24001) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19248) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12178) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4114) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25496) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14303) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17034) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15186) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28673) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15288) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2247) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20730) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20498) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17128) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10170) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13177) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23833) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25736) * $signed(input_fmap_34[7:0]) +
	( 5'sd 10) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19134) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8208) * $signed(input_fmap_40[7:0]) +
	( 11'sd 549) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5880) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4412) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31309) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3668) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25081) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2440) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4447) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24649) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12459) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29879) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8580) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2324) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24365) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21897) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5123) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25737) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10486) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31471) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7711) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6805) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25890) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7949) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12698) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8764) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20889) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10695) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21967) * $signed(input_fmap_89[7:0]) +
	( 9'sd 184) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4626) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14998) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20605) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28261) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5960) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1288) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23878) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32691) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31978) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13248) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10921) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24659) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1534) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18289) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25658) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21025) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3323) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9658) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3648) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32297) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16196) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26489) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6578) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19186) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17585) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31942) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 15'sd 9655) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14036) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23403) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1449) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5930) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10867) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17576) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13856) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3623) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9520) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30709) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22494) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28799) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19477) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29754) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30895) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29638) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10925) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21181) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5400) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31609) * $signed(input_fmap_34[7:0]) +
	( 10'sd 483) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24426) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6823) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11623) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1991) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10749) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7679) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25408) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10242) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11328) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20180) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20858) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1382) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18934) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_55[7:0]) +
	( 14'sd 8175) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1707) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5449) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12162) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31145) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28249) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31874) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16891) * $signed(input_fmap_67[7:0]) +
	( 11'sd 911) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15614) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15159) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14243) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11957) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11639) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1762) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5301) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8452) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22582) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31752) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9417) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4682) * $signed(input_fmap_90[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21697) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4403) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2978) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2130) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16284) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20936) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20202) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5793) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_102[7:0]) +
	( 9'sd 186) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8829) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22766) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12956) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12658) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26909) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17430) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32210) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7042) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8381) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11731) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12028) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27120) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17435) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7701) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10395) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31170) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10649) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 16'sd 24165) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22241) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4649) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11928) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3360) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23757) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23698) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32401) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16838) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1089) * $signed(input_fmap_12[7:0]) +
	( 11'sd 791) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28082) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4309) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18913) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30341) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28250) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26320) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23265) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3312) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12574) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32527) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8817) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7093) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8677) * $signed(input_fmap_38[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28722) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5775) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11326) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29866) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4845) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13572) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6874) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28722) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15109) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29188) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31300) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7732) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3936) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32622) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28181) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13574) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22970) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1160) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8807) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13481) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29109) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30364) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1867) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14475) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25154) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27405) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7401) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10410) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6348) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4982) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20987) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25151) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27663) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2845) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23349) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29996) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28329) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30786) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21814) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13336) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14117) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28181) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22659) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21961) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19839) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2144) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1365) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4193) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13394) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26507) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11440) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9481) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20381) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28543) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14026) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6150) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_123[7:0]) +
	( 14'sd 8089) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 16'sd 20469) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16481) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17580) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26234) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8638) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12770) * $signed(input_fmap_5[7:0]) +
	( 11'sd 695) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29098) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4960) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32731) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5001) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20901) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23165) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8521) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23931) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28108) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10068) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9069) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29492) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4491) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22726) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22865) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7816) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13372) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16717) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27869) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25077) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6216) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5142) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10303) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29921) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1602) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26742) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27852) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_53[7:0]) +
	( 11'sd 820) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6795) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7557) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26426) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8758) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29688) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11543) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3159) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23281) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22525) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_67[7:0]) +
	( 11'sd 653) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_69[7:0]) +
	( 9'sd 210) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9856) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14084) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22641) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5895) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12369) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23794) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20550) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17909) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5216) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23671) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6239) * $signed(input_fmap_86[7:0]) +
	( 10'sd 342) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26079) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23460) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27986) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28101) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11550) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32611) * $signed(input_fmap_100[7:0]) +
	( 11'sd 820) * $signed(input_fmap_101[7:0]) +
	( 11'sd 906) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10038) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5281) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22628) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29491) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21436) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18340) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20829) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19327) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18446) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18310) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22572) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7067) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4828) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27802) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18880) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20364) * $signed(input_fmap_123[7:0]) +
	( 9'sd 250) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1248) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 16'sd 22657) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30797) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4724) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2695) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21273) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28337) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3683) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1602) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6042) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31116) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13146) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4313) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28963) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18250) * $signed(input_fmap_28[7:0]) +
	( 10'sd 376) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3179) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10898) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26242) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6071) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7567) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9350) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20929) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11057) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6144) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26699) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18292) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12725) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20683) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1466) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1076) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12309) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27866) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3946) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24363) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8683) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28811) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20764) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19322) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31012) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20076) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15952) * $signed(input_fmap_83[7:0]) +
	( 13'sd 4055) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26542) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10996) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20158) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2425) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3985) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18676) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22068) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29052) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16154) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20007) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16077) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27926) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31337) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7591) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_113[7:0]) +
	( 11'sd 767) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28420) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12330) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1803) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9148) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28964) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24503) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10057) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 16'sd 30297) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11914) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26707) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30020) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19519) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1159) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2381) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5946) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17297) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22481) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23092) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14265) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20987) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16679) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7507) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11550) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13581) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26641) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10953) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17918) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5934) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24857) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29743) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1726) * $signed(input_fmap_39[7:0]) +
	( 11'sd 556) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7285) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28032) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27751) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31611) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2698) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4536) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4611) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15559) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30605) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29258) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32461) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28690) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3560) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18829) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7622) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9668) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32093) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31362) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7564) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13184) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_75[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27990) * $signed(input_fmap_77[7:0]) +
	( 10'sd 490) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14903) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3305) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29773) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16015) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27665) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8633) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29061) * $signed(input_fmap_91[7:0]) +
	( 12'sd 2037) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7045) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31452) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7474) * $signed(input_fmap_96[7:0]) +
	( 11'sd 768) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21215) * $signed(input_fmap_98[7:0]) +
	( 8'sd 122) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14418) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7696) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22188) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5355) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19063) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26279) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12174) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24867) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29686) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7775) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20876) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32542) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13762) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22926) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23798) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29166) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32138) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21708) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1336) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13821) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 16'sd 27581) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30497) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17384) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28738) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6039) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20446) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25240) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13361) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32706) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1711) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30334) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32048) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2429) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27509) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2285) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22981) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13977) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13528) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13861) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30874) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11390) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11508) * $signed(input_fmap_25[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3941) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13010) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20787) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8473) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18370) * $signed(input_fmap_34[7:0]) +
	( 14'sd 8058) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20359) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5698) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1265) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23996) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8485) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7223) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6167) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1355) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19588) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10004) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13631) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24040) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1561) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11493) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16992) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19305) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17008) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20486) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13637) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4225) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32680) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17424) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20941) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7475) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3510) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9305) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15657) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3807) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6315) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18145) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12354) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4405) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11788) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2255) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5847) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5226) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6113) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14128) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14484) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10587) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9238) * $signed(input_fmap_114[7:0]) +
	( 8'sd 92) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16210) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8743) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2755) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12614) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4449) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3104) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11573) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22132) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 11'sd 829) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5648) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9062) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24408) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18871) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6167) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26490) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16333) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30557) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22146) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15796) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8878) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15228) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12699) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23594) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14607) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28534) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22395) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26474) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10558) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22583) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32756) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17790) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13409) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22181) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7921) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26687) * $signed(input_fmap_37[7:0]) +
	( 11'sd 874) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31259) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17509) * $signed(input_fmap_40[7:0]) +
	( 11'sd 570) * $signed(input_fmap_41[7:0]) +
	( 14'sd 8032) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8262) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26789) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22285) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26051) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27787) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6350) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11823) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24399) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8865) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11403) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_63[7:0]) +
	( 4'sd 7) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5587) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32283) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30988) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2192) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2663) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18396) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1349) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17793) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20063) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12577) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26641) * $signed(input_fmap_82[7:0]) +
	( 11'sd 542) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29312) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6902) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4483) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13591) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26898) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13091) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10773) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25963) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8791) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22375) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8130) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21022) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31067) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17431) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21160) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15580) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2315) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7054) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9119) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11727) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28142) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5797) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2934) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18617) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18567) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9279) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30973) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28860) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14674) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21282) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24082) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15538) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 13'sd 4015) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13568) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25030) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28767) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13634) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11349) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28291) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7132) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12741) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18115) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15326) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7911) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1363) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28866) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_18[7:0]) +
	( 11'sd 738) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20832) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8791) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15344) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26658) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9779) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13750) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22774) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24742) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23835) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6376) * $signed(input_fmap_37[7:0]) +
	( 10'sd 416) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4503) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1993) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1082) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25555) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2788) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18838) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18832) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32646) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20784) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27023) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10641) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17558) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1687) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24512) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_61[7:0]) +
	( 11'sd 958) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14827) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32162) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22043) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23688) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6390) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26523) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12731) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22199) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22581) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10451) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11897) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16366) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5356) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16025) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30620) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_84[7:0]) +
	( 6'sd 20) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15646) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21552) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16697) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32289) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30769) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6641) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20963) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10837) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28916) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12172) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12551) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21079) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4573) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22724) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13487) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_112[7:0]) +
	( 4'sd 4) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17632) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28445) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11845) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10563) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30874) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18255) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22790) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17953) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 16'sd 28790) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4428) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3389) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17937) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30440) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17939) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25748) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17659) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13499) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26456) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15849) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18190) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10919) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30331) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20730) * $signed(input_fmap_21[7:0]) +
	( 11'sd 896) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2910) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15439) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12226) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21695) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8837) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19468) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8703) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27803) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17992) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16368) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9181) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12136) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27678) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2443) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21482) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9925) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2468) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10798) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15127) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23719) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9728) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12204) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20285) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22381) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19017) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9839) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4450) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30473) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15755) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29108) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27391) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23134) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13915) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5367) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9216) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1707) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19523) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6998) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9286) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1937) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1719) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8789) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4909) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26737) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24460) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5627) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1723) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1874) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21204) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8285) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26018) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32024) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5572) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23073) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_106[7:0]) +
	( 11'sd 649) * $signed(input_fmap_107[7:0]) +
	( 11'sd 563) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20836) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26985) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3012) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24073) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22525) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3556) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27736) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13936) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11906) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18999) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19367) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10434) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7711) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 16'sd 30688) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11990) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30399) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31870) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24903) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19476) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2452) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25593) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13460) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25960) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4600) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1100) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16207) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_22[7:0]) +
	( 11'sd 821) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25660) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27608) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5940) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9224) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4532) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4379) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7303) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31840) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27551) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7160) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19281) * $signed(input_fmap_36[7:0]) +
	( 11'sd 956) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28671) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16263) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18552) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5162) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23871) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4798) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22614) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19777) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22508) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2957) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1084) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17523) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23405) * $signed(input_fmap_56[7:0]) +
	( 11'sd 524) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22609) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17797) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2779) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_61[7:0]) +
	( 10'sd 313) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_63[7:0]) +
	( 11'sd 979) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22270) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1865) * $signed(input_fmap_66[7:0]) +
	( 10'sd 450) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26641) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18396) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22827) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21253) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_74[7:0]) +
	( 11'sd 794) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7240) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11203) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9427) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17811) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30620) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24252) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27967) * $signed(input_fmap_87[7:0]) +
	( 9'sd 205) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12243) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4232) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15882) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29613) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20513) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23617) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9006) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29144) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17388) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6777) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12024) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29926) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29454) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23999) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25848) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3071) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3563) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_121[7:0]) +
	( 10'sd 480) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25035) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24270) * $signed(input_fmap_125[7:0]) +
	( 11'sd 551) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 12'sd 1593) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32380) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_2[7:0]) +
	( 11'sd 751) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26820) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4747) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30011) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26329) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10842) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32039) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22002) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6151) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11928) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6386) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12366) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15747) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7027) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8488) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11192) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13847) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5448) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17867) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10629) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10094) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19477) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25250) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3865) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20475) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28813) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_40[7:0]) +
	( 10'sd 295) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5633) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23151) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18050) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14008) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28015) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27989) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25124) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15925) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4567) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_59[7:0]) +
	( 10'sd 257) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1691) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_65[7:0]) +
	( 10'sd 339) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23906) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11972) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21234) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6073) * $signed(input_fmap_70[7:0]) +
	( 9'sd 208) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14916) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26951) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29300) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29916) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14085) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32352) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25162) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21635) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3381) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13937) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24399) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3884) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27499) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28586) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9998) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15027) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12253) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7959) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21398) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20900) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20960) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19756) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22914) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2055) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18163) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29343) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11718) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9376) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4365) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10909) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19410) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13648) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22371) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 14'sd 7794) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27914) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10032) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31016) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17988) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3940) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12389) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30257) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1772) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27770) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30707) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30097) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7229) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4306) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26186) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23961) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17379) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20060) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24570) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16524) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21660) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25227) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19667) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29718) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2381) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19718) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18780) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8796) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16884) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3684) * $signed(input_fmap_45[7:0]) +
	( 14'sd 8075) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16172) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5938) * $signed(input_fmap_48[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15235) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10017) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8540) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31139) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30976) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27955) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6655) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10469) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5596) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26884) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16016) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20875) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29608) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13818) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11290) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30406) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28123) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6785) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3012) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28763) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24137) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6943) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13953) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24845) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3771) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12691) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11503) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16318) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1648) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10144) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5356) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21099) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19980) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3414) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19688) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29219) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21984) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4870) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25097) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22621) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17016) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8472) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26444) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3999) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_126[7:0]) +
	( 9'sd 196) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 16'sd 18879) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27489) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27989) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2215) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14921) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12975) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6626) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31165) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8907) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28271) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28727) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26852) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11676) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1574) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26749) * $signed(input_fmap_21[7:0]) +
	( 11'sd 870) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12893) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32532) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29955) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30384) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26312) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17159) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28904) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11951) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32316) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16466) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_39[7:0]) +
	( 10'sd 450) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6725) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17456) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13450) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13466) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2331) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8819) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21509) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9749) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12976) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19520) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5096) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32655) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27937) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7478) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23433) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18979) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15823) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17115) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6712) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29941) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1134) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31553) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30131) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31265) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20506) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4725) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31792) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8773) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19115) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23575) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8015) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27576) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8385) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32467) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16540) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4493) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5087) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8700) * $signed(input_fmap_98[7:0]) +
	( 11'sd 957) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19605) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14622) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31806) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20414) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30489) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20153) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18223) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24936) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23337) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27944) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3680) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6718) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15210) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11651) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15776) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30964) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 15'sd 8677) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26585) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20712) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_5[7:0]) +
	( 10'sd 299) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1047) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1143) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15116) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26175) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3624) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28504) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8710) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27001) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23786) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27870) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20552) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28366) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18639) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31824) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30418) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12179) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_33[7:0]) +
	( 11'sd 914) * $signed(input_fmap_34[7:0]) +
	( 14'sd 8167) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20805) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28556) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20171) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28561) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13091) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25305) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28856) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17256) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5687) * $signed(input_fmap_48[7:0]) +
	( 11'sd 755) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10252) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3694) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15296) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10850) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11131) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18710) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29661) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11741) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24576) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7031) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21703) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31753) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8718) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28795) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19732) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29286) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4367) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18641) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11664) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5814) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2772) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4340) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27095) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7942) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17125) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31632) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14163) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29340) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29500) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32333) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18436) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15980) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3073) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21480) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13389) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27226) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7095) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19428) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29527) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12455) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19992) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1786) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17201) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27731) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4354) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31249) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12969) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7277) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8927) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 16'sd 21735) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30423) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23900) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7125) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14650) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19222) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9266) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8523) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2752) * $signed(input_fmap_10[7:0]) +
	( 10'sd 412) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23919) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21464) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21905) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28161) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11137) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13354) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4276) * $signed(input_fmap_20[7:0]) +
	( 11'sd 526) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7783) * $signed(input_fmap_23[7:0]) +
	( 11'sd 514) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14699) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4766) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28978) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24996) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14480) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8934) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20195) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13677) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28536) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30137) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11914) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13071) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16165) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6822) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8379) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28853) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24026) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19999) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2747) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_50[7:0]) +
	( 7'sd 59) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16115) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4870) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23983) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28718) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27070) * $signed(input_fmap_58[7:0]) +
	( 10'sd 356) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11036) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25314) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18998) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3977) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26871) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8393) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17552) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11469) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5825) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1367) * $signed(input_fmap_79[7:0]) +
	( 10'sd 435) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26063) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10757) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3181) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31324) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6175) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2053) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9629) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23940) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2508) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15135) * $signed(input_fmap_92[7:0]) +
	( 10'sd 353) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25235) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13257) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29145) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1951) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21881) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5055) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31716) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13733) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18252) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24191) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5737) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29857) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30385) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23011) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19608) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19800) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15850) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3725) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22712) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28491) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19713) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 16'sd 23980) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30784) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30737) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8846) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6900) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28046) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10111) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8444) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22104) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21436) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30849) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26578) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31022) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32035) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21111) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5008) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10358) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18589) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25828) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5663) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14855) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17792) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26792) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6327) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23202) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24820) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13397) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5325) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23314) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9600) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13509) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12637) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17690) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31437) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15062) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7456) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29766) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8200) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4347) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27914) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11556) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11285) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31953) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30005) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3424) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16467) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3415) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12878) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5383) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6543) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23551) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11542) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32146) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9756) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15293) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2467) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24617) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15185) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19225) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22323) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21429) * $signed(input_fmap_90[7:0]) +
	( 11'sd 695) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20057) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19779) * $signed(input_fmap_94[7:0]) +
	( 6'sd 30) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25803) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16056) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19701) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25861) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7675) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3781) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15401) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25727) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27424) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8209) * $signed(input_fmap_116[7:0]) +
	( 11'sd 703) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11419) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19047) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8273) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32551) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20108) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5417) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 14'sd 7366) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_1[7:0]) +
	( 10'sd 500) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16114) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18835) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14070) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5188) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26178) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11228) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1961) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28834) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12845) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25798) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3187) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31878) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21718) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17087) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29260) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13993) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14836) * $signed(input_fmap_31[7:0]) +
	( 7'sd 50) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15412) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29165) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28398) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6243) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13646) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19316) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25396) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22645) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31252) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7527) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_52[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31186) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2720) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9745) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13709) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22387) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8459) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_61[7:0]) +
	( 11'sd 575) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14707) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30982) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23938) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20098) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23653) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13942) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29180) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17516) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11359) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6550) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13101) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26886) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32268) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8433) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9346) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_87[7:0]) +
	( 10'sd 366) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15330) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11071) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26226) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15037) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32416) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26892) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27071) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_98[7:0]) +
	( 11'sd 812) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19694) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3303) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26911) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6681) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23493) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14027) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2782) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1176) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14900) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27008) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11510) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6674) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24835) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31562) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6454) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24456) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19347) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25309) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11258) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9460) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12793) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 16'sd 26539) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20552) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27048) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31399) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23151) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16833) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21784) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10389) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32230) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16998) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30582) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18390) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27739) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15445) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1479) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_21[7:0]) +
	( 11'sd 677) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21648) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27430) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13238) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30004) * $signed(input_fmap_28[7:0]) +
	( 9'sd 253) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13547) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22605) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29219) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12056) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31335) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5458) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19577) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6438) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28666) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17965) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16167) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29736) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25803) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13569) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8597) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24740) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12074) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21932) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9217) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10205) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23430) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11423) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17758) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5963) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23324) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22242) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26881) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19882) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7296) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27426) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12769) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25343) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12535) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18688) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8662) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3789) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31279) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32166) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10829) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5847) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16070) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13199) * $signed(input_fmap_101[7:0]) +
	( 11'sd 993) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4583) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31694) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13883) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5408) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_109[7:0]) +
	( 11'sd 653) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_111[7:0]) +
	( 10'sd 441) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3431) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2140) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18581) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23150) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2412) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28292) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16063) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 15'sd 14117) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21533) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23194) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13657) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1976) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26259) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16497) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4916) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20688) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5365) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8852) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10395) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19727) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9043) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26788) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5491) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7973) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2602) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11594) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8760) * $signed(input_fmap_27[7:0]) +
	( 11'sd 745) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23392) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4683) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19241) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17490) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3678) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_35[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9167) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14353) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3290) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31896) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28509) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26099) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8961) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10624) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28761) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20926) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28715) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27997) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31038) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10241) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5204) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27594) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5881) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30754) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11548) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10828) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2221) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13432) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27693) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_77[7:0]) +
	( 11'sd 991) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24206) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28985) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_83[7:0]) +
	( 11'sd 1014) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24053) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27481) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19698) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7915) * $signed(input_fmap_88[7:0]) +
	( 11'sd 716) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21727) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24258) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9758) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5828) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13372) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6519) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28017) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22638) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6499) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21715) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23422) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17677) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12210) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_107[7:0]) +
	( 10'sd 421) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9800) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5516) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31460) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15085) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6847) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24101) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17232) * $signed(input_fmap_121[7:0]) +
	( 13'sd 4001) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9501) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26639) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12117) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 15'sd 11568) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18892) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5439) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30383) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22909) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13845) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8067) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23159) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31721) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18032) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1878) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13643) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16604) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5227) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30546) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29480) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18163) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7931) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18744) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13341) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29867) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12537) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2091) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13976) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10542) * $signed(input_fmap_39[7:0]) +
	( 9'sd 175) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13884) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23211) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23154) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3457) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14891) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5455) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28571) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23711) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13987) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13788) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2333) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17560) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29210) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26489) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11457) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14289) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25510) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4187) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22343) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12483) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13643) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5743) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_83[7:0]) +
	( 11'sd 811) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4667) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30905) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32515) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8468) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20673) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16712) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7464) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18603) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26754) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19664) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14656) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17729) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19401) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1578) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_104[7:0]) +
	( 9'sd 249) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5256) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16731) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19510) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20746) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16934) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5265) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13812) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17862) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8935) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16634) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_124[7:0]) +
	( 10'sd 265) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5590) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2548) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 16'sd 23953) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8197) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7098) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23330) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14776) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29673) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19095) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25446) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12420) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16559) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29573) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29231) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12635) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2408) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20664) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5219) * $signed(input_fmap_26[7:0]) +
	( 11'sd 833) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17701) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26767) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29787) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3141) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9921) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9804) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30716) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32513) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17576) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28078) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13697) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6930) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2311) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6320) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19893) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15533) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3340) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10922) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2666) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_61[7:0]) +
	( 11'sd 715) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1361) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26975) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26701) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3694) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23251) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_69[7:0]) +
	( 5'sd 11) * $signed(input_fmap_70[7:0]) +
	( 10'sd 437) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17900) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2440) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25501) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26593) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11012) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3278) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29561) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8846) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8832) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27499) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29809) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2770) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18640) * $signed(input_fmap_95[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27999) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28927) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31097) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14633) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23535) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23118) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16289) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31806) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20070) * $signed(input_fmap_110[7:0]) +
	( 10'sd 408) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28789) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17213) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24663) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5357) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7874) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7486) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9178) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25828) * $signed(input_fmap_122[7:0]) +
	( 11'sd 646) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3413) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11061) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2893) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 15'sd 10968) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5049) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23747) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12682) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16096) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21799) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3174) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_11[7:0]) +
	( 11'sd 572) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23402) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15040) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28064) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2474) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8909) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15715) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9573) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10057) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7475) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16035) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20578) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12640) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29584) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4645) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14152) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18013) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1267) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11994) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13518) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4915) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4752) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9581) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32070) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7570) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12305) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21697) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11914) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_51[7:0]) +
	( 12'sd 2046) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32476) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24763) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16489) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6627) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6253) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16314) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_64[7:0]) +
	( 13'sd 4046) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24100) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22158) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21870) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3230) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20089) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11164) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22632) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12052) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24351) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19813) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2426) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15070) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15560) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18745) * $signed(input_fmap_95[7:0]) +
	( 10'sd 452) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6697) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5742) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3847) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10864) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8420) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6045) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22725) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1453) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5636) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5221) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15436) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30807) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13782) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23003) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28425) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28245) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9811) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 11'sd 629) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31388) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5810) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30862) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20286) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8156) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_6[7:0]) +
	( 10'sd 355) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17864) * $signed(input_fmap_8[7:0]) +
	( 11'sd 870) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21431) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18087) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31051) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19342) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10437) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23132) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14990) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8668) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5018) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13311) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9291) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_25[7:0]) +
	( 9'sd 238) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13341) * $signed(input_fmap_28[7:0]) +
	( 10'sd 336) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31786) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31505) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5570) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32029) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32711) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10245) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15328) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29836) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5045) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19203) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29762) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23851) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9539) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16210) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16503) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2856) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19365) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29005) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12378) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19662) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19327) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26735) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15104) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9571) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17769) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24040) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8296) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25159) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20680) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17494) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2592) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18885) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6652) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13920) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15858) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16597) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16950) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26140) * $signed(input_fmap_91[7:0]) +
	( 13'sd 4030) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5243) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31890) * $signed(input_fmap_95[7:0]) +
	( 9'sd 204) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26325) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23231) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22026) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29400) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17551) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23654) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27017) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3734) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5773) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20863) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28327) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24083) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16501) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27647) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9267) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5579) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32418) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21986) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27356) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 16'sd 27571) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12904) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8347) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20865) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18349) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28929) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1832) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27187) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21808) * $signed(input_fmap_9[7:0]) +
	( 11'sd 846) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5845) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4625) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1181) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9034) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4638) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16925) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14665) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18908) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26314) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16253) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2670) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5878) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23541) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14811) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28835) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26291) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15560) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4699) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28532) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32445) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15561) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23319) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28108) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3117) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13486) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7722) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18233) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21744) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26418) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13394) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9710) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32349) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24223) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21021) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3948) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4372) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14659) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32380) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24663) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31054) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7622) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6242) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11761) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4683) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1924) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18561) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21506) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12584) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8723) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28096) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18680) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_94[7:0]) +
	( 7'sd 51) * $signed(input_fmap_95[7:0]) +
	( 11'sd 621) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2835) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26899) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20720) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5815) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3506) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8164) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15176) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11230) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6146) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20882) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2071) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20754) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22621) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27583) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21918) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22081) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25125) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16335) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24679) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28800) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31902) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6383) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27636) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_124[7:0]) +
	( 13'sd 4087) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26268) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15097) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 16'sd 23294) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28811) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13408) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4585) * $signed(input_fmap_3[7:0]) +
	( 9'sd 166) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25971) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27249) * $signed(input_fmap_6[7:0]) +
	( 11'sd 539) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16992) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20473) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7441) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20842) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_13[7:0]) +
	( 8'sd 114) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4687) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3748) * $signed(input_fmap_17[7:0]) +
	( 13'sd 4082) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22054) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10814) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6651) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2232) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1629) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29221) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25368) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16540) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26006) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30375) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5244) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13710) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15458) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15858) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32519) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22616) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12349) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19204) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32713) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22140) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17717) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1295) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29371) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26465) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4192) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2781) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6678) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15756) * $signed(input_fmap_57[7:0]) +
	( 11'sd 668) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12381) * $signed(input_fmap_59[7:0]) +
	( 10'sd 322) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_61[7:0]) +
	( 11'sd 593) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12915) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6837) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31553) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29196) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6185) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4297) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6257) * $signed(input_fmap_77[7:0]) +
	( 11'sd 597) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15805) * $signed(input_fmap_81[7:0]) +
	( 9'sd 128) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23711) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19645) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25670) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5507) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1117) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6669) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11042) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25689) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16518) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10994) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9612) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30135) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30051) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15295) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5398) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7644) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5188) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32147) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28742) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8208) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20650) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28674) * $signed(input_fmap_116[7:0]) +
	( 10'sd 462) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24726) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9915) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8270) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28507) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31742) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32690) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 16'sd 17721) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3644) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24746) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15110) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30084) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19846) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22888) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_11[7:0]) +
	( 11'sd 653) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19229) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22045) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5899) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11940) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5530) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25189) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27450) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19897) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28471) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16899) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19017) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29826) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30400) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9392) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27430) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15198) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_35[7:0]) +
	( 11'sd 558) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17035) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7022) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20626) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5829) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15335) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7344) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14672) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2244) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11358) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29942) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26751) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31236) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1107) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27846) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6760) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6267) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6561) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20378) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16838) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29045) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11084) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32453) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30200) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27171) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_72[7:0]) +
	( 9'sd 207) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31674) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3322) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27877) * $signed(input_fmap_78[7:0]) +
	( 10'sd 461) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9011) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21947) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28578) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28339) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25488) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_89[7:0]) +
	( 10'sd 451) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8754) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18704) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14336) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2469) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32543) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11340) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31854) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23150) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8919) * $signed(input_fmap_101[7:0]) +
	( 10'sd 291) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29498) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6888) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8136) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5478) * $signed(input_fmap_112[7:0]) +
	( 10'sd 509) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9180) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13189) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11936) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17271) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3018) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18027) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4330) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32586) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 16'sd 25512) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23842) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25204) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23190) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15593) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7130) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22456) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21374) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9392) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25343) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32540) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1739) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25591) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21740) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23154) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1264) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17945) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28079) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23701) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1409) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16664) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11724) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11032) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32267) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8688) * $signed(input_fmap_43[7:0]) +
	( 10'sd 388) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9625) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30229) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19973) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22505) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15781) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9703) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9045) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1238) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6861) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5906) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22121) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22029) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13883) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13558) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26340) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15010) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4788) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25563) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9349) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9055) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20789) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18604) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7364) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18393) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31667) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10146) * $signed(input_fmap_81[7:0]) +
	( 10'sd 346) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26954) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32446) * $signed(input_fmap_90[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18692) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2289) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17670) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30989) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3806) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3665) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30103) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22367) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28183) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2506) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14222) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4513) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29357) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9571) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3173) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24642) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27321) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14102) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12015) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29785) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1288) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 16'sd 31601) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29296) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4915) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_3[7:0]) +
	( 9'sd 143) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8094) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10766) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6319) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18123) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16947) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17006) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30470) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7824) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27243) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6987) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4491) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27274) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25272) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2555) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19584) * $signed(input_fmap_25[7:0]) +
	( 11'sd 983) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10497) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_28[7:0]) +
	( 11'sd 665) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21424) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31056) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28336) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29798) * $signed(input_fmap_35[7:0]) +
	( 11'sd 627) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3582) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2286) * $signed(input_fmap_38[7:0]) +
	( 11'sd 530) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26064) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25045) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30167) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12739) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32372) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10823) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29659) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5643) * $signed(input_fmap_49[7:0]) +
	( 10'sd 370) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3041) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1176) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28770) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5281) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25242) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11188) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31979) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18419) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21488) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4341) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28273) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6460) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6860) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11455) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1772) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6807) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31646) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21864) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12826) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12124) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24723) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2825) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9052) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16307) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30900) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2635) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14216) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9079) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10287) * $signed(input_fmap_103[7:0]) +
	( 11'sd 826) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19709) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25397) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5106) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_109[7:0]) +
	( 10'sd 287) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1045) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9640) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28198) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26228) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27303) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7038) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3771) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9044) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24089) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 15'sd 11927) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31463) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25368) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10138) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7646) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14210) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25194) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14750) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30010) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21777) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30074) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7870) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27866) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21383) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15451) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12529) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4609) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18495) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27253) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20440) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16306) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1442) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18633) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6541) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21022) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17435) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8008) * $signed(input_fmap_33[7:0]) +
	( 7'sd 35) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16868) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1536) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30380) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24032) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18182) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11880) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7937) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30591) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24362) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23584) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17713) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13327) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19078) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19576) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28775) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13835) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27047) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31568) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14171) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1931) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26226) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29075) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17745) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32597) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7425) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30131) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7200) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16406) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18037) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18363) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25101) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26119) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11110) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4549) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12597) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1266) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_87[7:0]) +
	( 10'sd 483) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31373) * $signed(input_fmap_89[7:0]) +
	( 10'sd 316) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25370) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29694) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13266) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18356) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18081) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_105[7:0]) +
	( 11'sd 559) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7800) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30571) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12344) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5266) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29408) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16698) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10748) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31316) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1952) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8230) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 16'sd 18774) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24059) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28049) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9157) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25633) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5411) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12116) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30849) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23125) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14369) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_20[7:0]) +
	( 11'sd 638) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13798) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7854) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3838) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8452) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15396) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10396) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22471) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24122) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30773) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4769) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16916) * $signed(input_fmap_37[7:0]) +
	( 11'sd 818) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4776) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_40[7:0]) +
	( 11'sd 1007) * $signed(input_fmap_41[7:0]) +
	( 6'sd 20) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18284) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18566) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5678) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13412) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11225) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24842) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2421) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18265) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27094) * $signed(input_fmap_54[7:0]) +
	( 7'sd 33) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8709) * $signed(input_fmap_56[7:0]) +
	( 9'sd 152) * $signed(input_fmap_57[7:0]) +
	( 10'sd 332) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19807) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8493) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1955) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20152) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14560) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10224) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26179) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19136) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14588) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1052) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10422) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29917) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8097) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9198) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13012) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3708) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12566) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13114) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16349) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21638) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2442) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29232) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16513) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7765) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5186) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11988) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31225) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17499) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30592) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29661) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13674) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22259) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16343) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25925) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27269) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17051) * $signed(input_fmap_119[7:0]) +
	( 11'sd 950) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15879) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26388) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23807) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_125[7:0]) +
	( 15'sd 16169) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18239) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 15'sd 14855) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_2[7:0]) +
	( 11'sd 900) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3553) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3013) * $signed(input_fmap_7[7:0]) +
	( 11'sd 512) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24533) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22565) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24728) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14337) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21300) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16048) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3182) * $signed(input_fmap_20[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6599) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7868) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13313) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29987) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19285) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19305) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2774) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12174) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16410) * $signed(input_fmap_38[7:0]) +
	( 7'sd 46) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24726) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8439) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9467) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32440) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16398) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_49[7:0]) +
	( 11'sd 611) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21831) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12563) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18734) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14237) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20192) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15952) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24707) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23751) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9871) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9120) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26628) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24948) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10787) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10433) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32157) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31138) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19672) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28372) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17789) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15335) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7568) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30042) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29561) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3161) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8600) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25611) * $signed(input_fmap_91[7:0]) +
	( 8'sd 100) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29180) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27283) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9587) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19778) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30072) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10995) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29279) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23071) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29823) * $signed(input_fmap_107[7:0]) +
	( 8'sd 122) * $signed(input_fmap_108[7:0]) +
	( 10'sd 496) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11442) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11426) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14770) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15976) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22809) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7431) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2723) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27090) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 16'sd 31067) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4781) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14447) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26631) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5943) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21505) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4385) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16149) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13485) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15364) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21711) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1574) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31412) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28245) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9895) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20842) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20992) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23915) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26064) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1670) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8542) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22165) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20473) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9572) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4149) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20753) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23451) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12190) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13884) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14452) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13187) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29256) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3421) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25236) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23799) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18369) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16919) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25784) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25034) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16590) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18416) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5566) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9870) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21188) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31285) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15825) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11865) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23481) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13439) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13202) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25495) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5124) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9704) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24513) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10188) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8707) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9410) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26332) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4946) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12478) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30951) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27784) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15791) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3619) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31798) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4875) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15915) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_111[7:0]) +
	( 9'sd 248) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20681) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27163) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9278) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3310) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1829) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3062) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16458) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24875) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 15'sd 16100) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15245) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16724) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29505) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16909) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28986) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20779) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9000) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10018) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30369) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28358) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6029) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14598) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26410) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3217) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22297) * $signed(input_fmap_20[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9663) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19712) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18605) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14351) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1043) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19697) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18766) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23526) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30406) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16804) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13635) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32223) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26969) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25454) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29284) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1887) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25716) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23970) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23190) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8842) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6577) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16307) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22533) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32449) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11013) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28059) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27617) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19507) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19556) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25043) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9068) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29133) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2153) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32720) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9544) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15970) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19190) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20271) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11545) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8582) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10577) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16536) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2817) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28023) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31842) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29811) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29217) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28308) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27019) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29073) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6448) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20667) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2788) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25545) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8167) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2071) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12082) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31199) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24406) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32201) * $signed(input_fmap_119[7:0]) +
	( 9'sd 136) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11686) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15709) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 16'sd 30323) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9211) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25660) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17864) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31892) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9393) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30910) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24415) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_16[7:0]) +
	( 11'sd 897) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19440) * $signed(input_fmap_18[7:0]) +
	( 12'sd 2032) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31830) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7849) * $signed(input_fmap_22[7:0]) +
	( 10'sd 353) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30033) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28597) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16937) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25369) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11722) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29508) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4905) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23829) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6313) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31979) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6190) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28092) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24001) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_40[7:0]) +
	( 14'sd 8040) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7662) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13062) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22446) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16053) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15094) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13637) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16762) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13041) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21619) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3572) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27577) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14761) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27510) * $signed(input_fmap_58[7:0]) +
	( 11'sd 658) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9598) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28448) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28136) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27636) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13518) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26304) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22372) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23150) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26015) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14904) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26623) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15161) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24765) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25809) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3827) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22127) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25223) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3776) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9760) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20707) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8096) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23743) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12121) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29064) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13422) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7435) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26179) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9606) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23396) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25098) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27738) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17421) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26970) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6917) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4210) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12891) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_110[7:0]) +
	( 11'sd 753) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9068) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32450) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14679) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20246) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15134) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20452) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18563) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17845) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4611) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 16'sd 24987) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11244) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17400) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_11[7:0]) +
	( 10'sd 268) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3651) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17666) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7425) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3258) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24191) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3042) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26296) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14555) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28765) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13804) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22334) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32280) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16023) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20506) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26434) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4965) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18158) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20056) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26204) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22325) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_47[7:0]) +
	( 11'sd 984) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15265) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28562) * $signed(input_fmap_51[7:0]) +
	( 11'sd 861) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19954) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30987) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18736) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26083) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22276) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31959) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28700) * $signed(input_fmap_66[7:0]) +
	( 10'sd 393) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_69[7:0]) +
	( 11'sd 795) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21148) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30762) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19898) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30397) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5948) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19795) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12846) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28224) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20140) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26711) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20818) * $signed(input_fmap_87[7:0]) +
	( 9'sd 176) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21256) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24150) * $signed(input_fmap_91[7:0]) +
	( 11'sd 970) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6818) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28412) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6615) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22795) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16627) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_101[7:0]) +
	( 9'sd 220) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6646) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29312) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14853) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2975) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7715) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27231) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1498) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19959) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14980) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16681) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 16'sd 23475) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22166) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8465) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29581) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5921) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6485) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24265) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9671) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15039) * $signed(input_fmap_10[7:0]) +
	( 7'sd 35) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_12[7:0]) +
	( 13'sd 4086) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1307) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10336) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26986) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12365) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12848) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30629) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3884) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30126) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4738) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5916) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24219) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32225) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24543) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28444) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21742) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18950) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12424) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19170) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24714) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1689) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28617) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10736) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8860) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16906) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17859) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14556) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31181) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3360) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16067) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9911) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28806) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24324) * $signed(input_fmap_64[7:0]) +
	( 11'sd 711) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19403) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17832) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19227) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24956) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31401) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16181) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11420) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14686) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10721) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20084) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18529) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4983) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17439) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6745) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12870) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1846) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15137) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9075) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9741) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11736) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15957) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23047) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1143) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1644) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27855) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28517) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19196) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18706) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32484) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11240) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17567) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14459) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3598) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7531) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15951) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31226) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25404) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22722) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11244) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16037) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5659) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25514) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15224) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22657) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12157) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29285) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12456) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 13'sd 2854) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30734) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17856) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13090) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24127) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20102) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_10[7:0]) +
	( 11'sd 831) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4852) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31027) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32317) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28157) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31217) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2955) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24428) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31264) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11753) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11554) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2199) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16762) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11090) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19834) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3857) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7565) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13507) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31289) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13225) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32243) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23458) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27421) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7161) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22616) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23469) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26224) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25082) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28452) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11888) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20235) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1977) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8410) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28416) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32273) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31841) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13300) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18263) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3437) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20779) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18258) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4290) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27940) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9264) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18713) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8370) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25389) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24275) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27670) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13640) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14036) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1577) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30993) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13007) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9842) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4313) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11108) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24339) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7530) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15159) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25694) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8524) * $signed(input_fmap_101[7:0]) +
	( 10'sd 416) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29131) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2510) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12439) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29455) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22828) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12423) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30018) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8053) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13634) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28964) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18238) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31397) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11060) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26806) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22348) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31179) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2687) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32575) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 15'sd 8490) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26229) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12735) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23112) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7694) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25719) * $signed(input_fmap_10[7:0]) +
	( 7'sd 37) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1989) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9030) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19733) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25180) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1148) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17662) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28576) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1480) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26388) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_31[7:0]) +
	( 9'sd 134) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30882) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24008) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27757) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3573) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21318) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27691) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18603) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9619) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9537) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21043) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28373) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20291) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27177) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11829) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2755) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1064) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10012) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19397) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9296) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16358) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23968) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25448) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12400) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18068) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9145) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1593) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12236) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12369) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20357) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30796) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18357) * $signed(input_fmap_84[7:0]) +
	( 11'sd 560) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16326) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11458) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9950) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28304) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25258) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24085) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14314) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1616) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29280) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10821) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8667) * $signed(input_fmap_100[7:0]) +
	( 11'sd 752) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1220) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22682) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26506) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18196) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32389) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28650) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18308) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11881) * $signed(input_fmap_115[7:0]) +
	( 13'sd 4048) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17527) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16280) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11725) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22153) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26254) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17633) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 15'sd 12087) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16165) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32564) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16702) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18552) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7176) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27991) * $signed(input_fmap_13[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21741) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13281) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17743) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6066) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31419) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18485) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26770) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21434) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9158) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26184) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23738) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16335) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7591) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25344) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9012) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26800) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16660) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2822) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16320) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30538) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22252) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10565) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32460) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18202) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11995) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21532) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15441) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25848) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24384) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17516) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18299) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20340) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16695) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13109) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7355) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31580) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5380) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24525) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18368) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26977) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4512) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8795) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1144) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20228) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6848) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30168) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27072) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15121) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2462) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14732) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21577) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4149) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_96[7:0]) +
	( 10'sd 498) * $signed(input_fmap_97[7:0]) +
	( 11'sd 656) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8617) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13885) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6102) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8805) * $signed(input_fmap_104[7:0]) +
	( 7'sd 53) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32280) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1249) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8335) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_114[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_116[7:0]) +
	( 10'sd 336) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32668) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27795) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11258) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23418) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17372) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30387) * $signed(input_fmap_126[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 13'sd 3801) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27348) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16368) * $signed(input_fmap_4[7:0]) +
	( 11'sd 949) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17467) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27266) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21143) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29214) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15657) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7445) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11505) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24226) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1955) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_20[7:0]) +
	( 11'sd 538) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20173) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20940) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_27[7:0]) +
	( 10'sd 403) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27933) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12357) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5058) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29427) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2256) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31382) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25028) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13854) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15906) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4856) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21473) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26815) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30122) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23576) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18509) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14431) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11555) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17046) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2147) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7522) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15813) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23268) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15508) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19190) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19557) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19172) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27387) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8994) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4377) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_77[7:0]) +
	( 11'sd 552) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8060) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26250) * $signed(input_fmap_81[7:0]) +
	( 11'sd 996) * $signed(input_fmap_82[7:0]) +
	( 11'sd 574) * $signed(input_fmap_83[7:0]) +
	( 11'sd 793) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6599) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16774) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25927) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26565) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24641) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17578) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29521) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6642) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20424) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31238) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21028) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31349) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6996) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_102[7:0]) +
	( 13'sd 4058) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6213) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30221) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2602) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21599) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16138) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31561) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11040) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14947) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25908) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30131) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13570) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_121[7:0]) +
	( 10'sd 272) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18561) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9142) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27845) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31534) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 15'sd 9422) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17642) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13882) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19229) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13895) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19245) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12291) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20369) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2126) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23435) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10719) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17473) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2454) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19929) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18462) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15474) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5808) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21400) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13884) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15625) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8424) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15939) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24884) * $signed(input_fmap_33[7:0]) +
	( 11'sd 774) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10553) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1871) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4781) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19425) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16695) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20185) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31391) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5355) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5526) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32730) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5810) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30793) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26926) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27499) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12213) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5299) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1664) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8606) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22721) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15353) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15265) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_68[7:0]) +
	( 11'sd 991) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2632) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16927) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17863) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13134) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17416) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7078) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1591) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11387) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31833) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5300) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25345) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29134) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26542) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9045) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32509) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30865) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7902) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17965) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11672) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24618) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21134) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24306) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10673) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31595) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5408) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30190) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9860) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30919) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26278) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14543) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9950) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6276) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25169) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12239) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4706) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13806) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_121[7:0]) +
	( 13'sd 4090) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31776) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13560) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 7'sd 46) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31137) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29325) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5440) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9537) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15377) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7191) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5220) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7788) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16691) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7736) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1282) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18612) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2579) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12998) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11537) * $signed(input_fmap_20[7:0]) +
	( 10'sd 256) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3184) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4489) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28271) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15081) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27740) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8902) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11884) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31661) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26135) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32343) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24403) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31662) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26037) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11916) * $signed(input_fmap_48[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24739) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30713) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19477) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14124) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13601) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24289) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20177) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29682) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31589) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16573) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17587) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20757) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20237) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32719) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15710) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12835) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9962) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14115) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24391) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20301) * $signed(input_fmap_81[7:0]) +
	( 11'sd 519) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13803) * $signed(input_fmap_84[7:0]) +
	( 11'sd 595) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29206) * $signed(input_fmap_86[7:0]) +
	( 9'sd 253) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29330) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29144) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26941) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11186) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13041) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11536) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16510) * $signed(input_fmap_94[7:0]) +
	( 11'sd 883) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14742) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21402) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16388) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1081) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20254) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13216) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26120) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5207) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10078) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23562) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8921) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20670) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10510) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14776) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5052) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13095) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 15'sd 10089) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24861) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27707) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5284) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29400) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23796) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16165) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_10[7:0]) +
	( 11'sd 590) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2638) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13533) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1279) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4151) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18405) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22082) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19563) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25248) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20116) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7566) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19224) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10529) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14940) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24537) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8738) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20615) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23377) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14899) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14632) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2596) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6281) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19125) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26511) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20049) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11865) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25574) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11969) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23952) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21717) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31450) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5685) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25157) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18042) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8014) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26126) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23513) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28032) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2820) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30556) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12821) * $signed(input_fmap_68[7:0]) +
	( 11'sd 535) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7588) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30553) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18887) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6478) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12404) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25737) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28127) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28657) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14680) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9700) * $signed(input_fmap_90[7:0]) +
	( 14'sd 8086) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13713) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4226) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14270) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26097) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23316) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22232) * $signed(input_fmap_101[7:0]) +
	( 11'sd 537) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18356) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16518) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28032) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14416) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_107[7:0]) +
	( 11'sd 734) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17005) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15853) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20374) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6756) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19296) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12770) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12998) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11322) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17675) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30460) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11732) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 16'sd 30503) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4949) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28472) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24321) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21272) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26327) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21079) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18519) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27278) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10819) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31910) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30872) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18995) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30125) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26636) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21462) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16657) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23319) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27830) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19907) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2283) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8890) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29062) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10767) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14443) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31780) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24850) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9921) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20138) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2255) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10558) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24811) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4878) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31463) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17314) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9088) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13245) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29055) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18190) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10716) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13402) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28972) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7449) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7185) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12686) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32243) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16611) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4464) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26528) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31822) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13305) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19429) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25733) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2928) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20574) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15437) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1466) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30391) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14137) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32303) * $signed(input_fmap_88[7:0]) +
	( 11'sd 1013) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31532) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21663) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28759) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17937) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_96[7:0]) +
	( 11'sd 802) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14429) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10977) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25563) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28286) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9921) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2713) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22887) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10317) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_107[7:0]) +
	( 11'sd 796) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17102) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18182) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27982) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27861) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7725) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30902) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17651) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29377) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27154) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1578) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14560) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22263) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31593) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10911) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11586) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28124) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16654) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 16'sd 30464) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29327) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19504) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14733) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18030) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5492) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28930) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_11[7:0]) +
	( 11'sd 588) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25121) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18683) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28339) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26794) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32464) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15264) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16972) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18162) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23361) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4119) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7687) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17640) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18091) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19546) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6201) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16878) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12580) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28892) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9022) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13993) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5593) * $signed(input_fmap_41[7:0]) +
	( 10'sd 426) * $signed(input_fmap_42[7:0]) +
	( 11'sd 822) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31276) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16087) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6923) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2300) * $signed(input_fmap_49[7:0]) +
	( 8'sd 95) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12987) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23300) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31326) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24077) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22910) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24030) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18380) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22813) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16761) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23751) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31685) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1659) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16383) * $signed(input_fmap_67[7:0]) +
	( 11'sd 650) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25339) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7558) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3447) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12677) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13993) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4403) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8405) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20661) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9964) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7788) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12879) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29345) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28127) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_93[7:0]) +
	( 11'sd 547) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25387) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27448) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7910) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4464) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12974) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25822) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23315) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17304) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28451) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32241) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10876) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22504) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3039) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9727) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27104) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7218) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3401) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17833) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29134) * $signed(input_fmap_125[7:0]) +
	( 11'sd 518) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2317) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 14'sd 7825) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8701) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19830) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_5[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32573) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6112) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5756) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8801) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23191) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12094) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23568) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11834) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23341) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15591) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18201) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2677) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32464) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23423) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1642) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9642) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6214) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5294) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11471) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32760) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7921) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13526) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12777) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3588) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2971) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14354) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25533) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19918) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32708) * $signed(input_fmap_53[7:0]) +
	( 11'sd 1004) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14182) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23100) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22775) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19671) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5645) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2676) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12502) * $signed(input_fmap_65[7:0]) +
	( 11'sd 717) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2808) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24176) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23321) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4578) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32464) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16134) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24440) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5622) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6766) * $signed(input_fmap_80[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9961) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15434) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2861) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30775) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30242) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27421) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28099) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1228) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5261) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9500) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3416) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17387) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17410) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17798) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14192) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2694) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5170) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9977) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22662) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15961) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30098) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18818) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13579) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26466) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 16'sd 31281) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26906) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7612) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23585) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3920) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5112) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24981) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31787) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20203) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15082) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11654) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25140) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18351) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9886) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20780) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29369) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6020) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24646) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15877) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4193) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19802) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11128) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16430) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27891) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11529) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11005) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22685) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19547) * $signed(input_fmap_44[7:0]) +
	( 11'sd 679) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10818) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10776) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15708) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14309) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18280) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23095) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21545) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1811) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26288) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6421) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2501) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16876) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11020) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15016) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32425) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10331) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20437) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16320) * $signed(input_fmap_70[7:0]) +
	( 9'sd 142) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24467) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19083) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12753) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32430) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19828) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19669) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14462) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18101) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13828) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17120) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22298) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_97[7:0]) +
	( 11'sd 690) * $signed(input_fmap_98[7:0]) +
	( 9'sd 218) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18236) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3255) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19322) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2805) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22015) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17646) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20529) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22906) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28966) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8176) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2986) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19931) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23018) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25461) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4144) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8620) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25352) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16732) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25050) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 11'sd 739) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7434) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30925) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13649) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9881) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2373) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15649) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2885) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17691) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28296) * $signed(input_fmap_16[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26010) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18612) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19360) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15106) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19861) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18347) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16056) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31789) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16288) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21578) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3801) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_37[7:0]) +
	( 11'sd 614) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12366) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14036) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24109) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5171) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5816) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1621) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11472) * $signed(input_fmap_47[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16223) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4756) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25345) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5537) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30452) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32550) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21573) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23582) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18873) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_59[7:0]) +
	( 10'sd 459) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29368) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5610) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5875) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10713) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8008) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1040) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17122) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_76[7:0]) +
	( 11'sd 750) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13964) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16294) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30590) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1280) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5421) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22859) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12461) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7956) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23992) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26723) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15642) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19402) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8836) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31477) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9718) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26326) * $signed(input_fmap_100[7:0]) +
	( 9'sd 223) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27865) * $signed(input_fmap_102[7:0]) +
	( 9'sd 247) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7459) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21962) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17744) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31125) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10605) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24463) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20375) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31364) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22469) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1122) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10995) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28478) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4775) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 11'sd 708) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14385) * $signed(input_fmap_1[7:0]) +
	( 11'sd 714) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17780) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32719) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15867) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8970) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13341) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28762) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4561) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18405) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18465) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_20[7:0]) +
	( 11'sd 813) * $signed(input_fmap_21[7:0]) +
	( 11'sd 748) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13825) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10988) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19506) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17232) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13658) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7158) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12158) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26882) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_35[7:0]) +
	( 10'sd 437) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9079) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27916) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22450) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30930) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25930) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9707) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5461) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2462) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7750) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18839) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17739) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24232) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1590) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7009) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8141) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6472) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11027) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6310) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9020) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8607) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20274) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21254) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16257) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31913) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19520) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2673) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28647) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31739) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14583) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28177) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11572) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18219) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25696) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11374) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21808) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22717) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19373) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21306) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14930) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28695) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10367) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20946) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9536) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1707) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7298) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9930) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18075) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19850) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25984) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30566) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20649) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9508) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13785) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24989) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30176) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 11'sd 759) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_1[7:0]) +
	( 10'sd 488) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24662) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7914) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19088) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4984) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29892) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18239) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_14[7:0]) +
	( 10'sd 274) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3544) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10303) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30662) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23327) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17179) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14181) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13918) * $signed(input_fmap_28[7:0]) +
	( 11'sd 940) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6095) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13281) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5019) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32690) * $signed(input_fmap_34[7:0]) +
	( 11'sd 996) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5079) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30917) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17231) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11650) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26717) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26763) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4719) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29980) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20612) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9891) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31700) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25508) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25344) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1129) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3171) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4815) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11204) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27877) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25586) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20807) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29367) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13744) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9559) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9515) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28188) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32268) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10140) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26880) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1143) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12588) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8469) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5804) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13089) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7431) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32708) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21244) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10123) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15987) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5036) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10085) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21415) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23597) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23000) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27056) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20127) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22302) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1693) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7239) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24573) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26490) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26004) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30508) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8283) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28220) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15270) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2174) * $signed(input_fmap_125[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_126[7:0]) +
	( 11'sd 978) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 16'sd 28337) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29030) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30777) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_3[7:0]) +
	( 10'sd 427) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1215) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27263) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6707) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17969) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13282) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32521) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10242) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23451) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3963) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29167) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13954) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27935) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14884) * $signed(input_fmap_30[7:0]) +
	( 11'sd 730) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17956) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22887) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28378) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13669) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8306) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21248) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2936) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28795) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20341) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7826) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26751) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21744) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_51[7:0]) +
	( 10'sd 451) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9206) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18244) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17593) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25841) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9839) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24223) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2582) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27739) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7464) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6555) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_67[7:0]) +
	( 9'sd 164) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13814) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27377) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2947) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22474) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14067) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25112) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11775) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10832) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30793) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10744) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9250) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22119) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_91[7:0]) +
	( 9'sd 181) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22419) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12179) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21909) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28286) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19558) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7325) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14402) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15882) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23371) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3335) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5546) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20923) * $signed(input_fmap_109[7:0]) +
	( 11'sd 565) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28188) * $signed(input_fmap_111[7:0]) +
	( 11'sd 622) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16395) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19716) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17057) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22955) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1974) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1416) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19465) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17622) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 16'sd 22515) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9253) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26321) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6800) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26174) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5664) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15996) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18049) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1769) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1474) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2630) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30808) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4347) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26287) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21032) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10358) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23439) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29105) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28033) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7633) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1974) * $signed(input_fmap_27[7:0]) +
	( 11'sd 592) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32436) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23393) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7387) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22266) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24388) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10559) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21546) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9731) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2647) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4716) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28207) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23656) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5563) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4431) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1875) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1203) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17920) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7370) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3651) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21885) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12751) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10357) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10124) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7922) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27740) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31057) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7168) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22129) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27467) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4687) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23440) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16716) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1233) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7611) * $signed(input_fmap_91[7:0]) +
	( 9'sd 239) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26712) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20396) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7445) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6620) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27140) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23139) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21895) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14819) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4618) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_111[7:0]) +
	( 10'sd 308) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31237) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32294) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7080) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23107) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7541) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19912) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10012) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29131) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23814) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25538) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 15'sd 12656) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19484) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22082) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21479) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12261) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14226) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9626) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2402) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31061) * $signed(input_fmap_12[7:0]) +
	( 7'sd 63) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31093) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8361) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23006) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8439) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29659) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8276) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8014) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29311) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14096) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28499) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12206) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32560) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24858) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32301) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24984) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18659) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7589) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7584) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16586) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3132) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13168) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21843) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4429) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25427) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29892) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11475) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14066) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8858) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6314) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18295) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24375) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31149) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11157) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23895) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23100) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9771) * $signed(input_fmap_63[7:0]) +
	( 10'sd 372) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15374) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32156) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13261) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13940) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13899) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16960) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11348) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10388) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30694) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14661) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13529) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11693) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3907) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1642) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11192) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9846) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11266) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1484) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9137) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7141) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22107) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17680) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4342) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27837) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27919) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9467) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17184) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3478) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4208) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13114) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6177) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23576) * $signed(input_fmap_116[7:0]) +
	( 11'sd 878) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_119[7:0]) +
	( 10'sd 343) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19361) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31607) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31764) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23419) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19444) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 16'sd 22981) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15633) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13262) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24827) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30727) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4195) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23516) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19436) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32376) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8500) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13177) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5703) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28890) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21141) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7372) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10012) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19563) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19470) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26211) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15609) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24615) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23672) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29567) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31478) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_38[7:0]) +
	( 9'sd 197) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13769) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20143) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31942) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32211) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30558) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24285) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23310) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2497) * $signed(input_fmap_50[7:0]) +
	( 8'sd 96) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24892) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13939) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28795) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11389) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32172) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16749) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16188) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24598) * $signed(input_fmap_72[7:0]) +
	( 11'sd 758) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20150) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17511) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4140) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9017) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18273) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10076) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32593) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7198) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15302) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13664) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7844) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11945) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13385) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23902) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32616) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23274) * $signed(input_fmap_102[7:0]) +
	( 10'sd 276) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20680) * $signed(input_fmap_105[7:0]) +
	( 10'sd 383) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32400) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3941) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27011) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21747) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_114[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15542) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9177) * $signed(input_fmap_117[7:0]) +
	( 9'sd 237) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21202) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24650) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23822) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11263) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29625) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 16'sd 28670) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26566) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27048) * $signed(input_fmap_4[7:0]) +
	( 11'sd 781) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27228) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5794) * $signed(input_fmap_7[7:0]) +
	( 9'sd 195) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8581) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6371) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18448) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11258) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23602) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9286) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17480) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10355) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3612) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27134) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22471) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11505) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_31[7:0]) +
	( 11'sd 556) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5743) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12639) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12652) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26693) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18116) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24872) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14097) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17713) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23954) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28482) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_52[7:0]) +
	( 9'sd 175) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9281) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18604) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12648) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30288) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17674) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4283) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11257) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4918) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21786) * $signed(input_fmap_66[7:0]) +
	( 11'sd 812) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23255) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30546) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25576) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9987) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19591) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21594) * $signed(input_fmap_74[7:0]) +
	( 10'sd 458) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32699) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13383) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28536) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4959) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21539) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25733) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18180) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11424) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_88[7:0]) +
	( 9'sd 201) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4249) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29638) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7127) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_93[7:0]) +
	( 10'sd 332) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12382) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4360) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14857) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15268) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11873) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4563) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18749) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1884) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24984) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2393) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2392) * $signed(input_fmap_106[7:0]) +
	( 11'sd 905) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7824) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13858) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31697) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27656) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12257) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14453) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18671) * $signed(input_fmap_120[7:0]) +
	( 13'sd 4002) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29121) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15096) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28529) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16388) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 16'sd 23213) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3808) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3348) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4398) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24486) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3686) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17045) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29515) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5785) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7743) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11973) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17114) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3598) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19628) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7618) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29642) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1701) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14965) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30123) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9893) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3486) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23867) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10177) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8508) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8619) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23942) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20080) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15749) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4813) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30730) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27074) * $signed(input_fmap_46[7:0]) +
	( 11'sd 549) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1978) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14372) * $signed(input_fmap_53[7:0]) +
	( 10'sd 349) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16970) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27154) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5946) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27506) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13628) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10394) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5876) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_65[7:0]) +
	( 11'sd 642) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16929) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27671) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22759) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21547) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5164) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3650) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11079) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32278) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22634) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7265) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30705) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27881) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16051) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26024) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9687) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23501) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21658) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19337) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24858) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_100[7:0]) +
	( 11'sd 586) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12253) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11086) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30003) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12463) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14561) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32710) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5846) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22167) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12354) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16986) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29343) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10914) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7016) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28827) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31232) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23668) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22767) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24779) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4700) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 14'sd 7713) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23953) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26297) * $signed(input_fmap_2[7:0]) +
	( 10'sd 269) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9418) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9497) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22789) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9012) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10580) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26653) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28906) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2795) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9638) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16011) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11251) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13418) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12939) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8841) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29040) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2160) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9142) * $signed(input_fmap_33[7:0]) +
	( 9'sd 244) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2141) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4399) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26233) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7935) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26413) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18294) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_48[7:0]) +
	( 10'sd 385) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25750) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28563) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12662) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22008) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19201) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12279) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30777) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26336) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1991) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10643) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24776) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17250) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29792) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4387) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_72[7:0]) +
	( 11'sd 784) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2387) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5670) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3251) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32258) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19157) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7644) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13417) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26957) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9672) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21492) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10828) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18588) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7995) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13435) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29379) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10577) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7755) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14255) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17902) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20070) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25727) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32733) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6754) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13700) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7723) * $signed(input_fmap_106[7:0]) +
	( 10'sd 434) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2863) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26094) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20881) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17082) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30278) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6340) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2501) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16128) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3828) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22452) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29059) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15144) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 16'sd 26863) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12160) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10751) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20286) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8415) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28342) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16597) * $signed(input_fmap_9[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3634) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13496) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_14[7:0]) +
	( 10'sd 382) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5886) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28329) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15392) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13055) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26762) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23271) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18121) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11553) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_27[7:0]) +
	( 9'sd 242) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14609) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5294) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10085) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2342) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27690) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25932) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15278) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31417) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24698) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20124) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7509) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11885) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12091) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28630) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12097) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29944) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29215) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8772) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24769) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6371) * $signed(input_fmap_71[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12673) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29062) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18531) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22113) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5416) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29860) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2859) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21575) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27006) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21829) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1307) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13502) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25017) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18414) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21448) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2856) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2827) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27704) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26983) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28876) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_102[7:0]) +
	( 11'sd 654) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18252) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16117) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24889) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26968) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15021) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28414) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24194) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12807) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32718) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13189) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23329) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16730) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16843) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30119) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22086) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15273) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2092) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 14'sd 6016) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7321) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9297) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7394) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12786) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16008) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16312) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28059) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7863) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17586) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27356) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23734) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3224) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4530) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23421) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8570) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1657) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27580) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24299) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25630) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30124) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31448) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31094) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6608) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17585) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14474) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30876) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18556) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31710) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7403) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14351) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29417) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6372) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_56[7:0]) +
	( 11'sd 605) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8859) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20903) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17121) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21931) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14892) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18390) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30888) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27264) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_71[7:0]) +
	( 8'sd 114) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21757) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14266) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6821) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15263) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9340) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29347) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13057) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20615) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31240) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3991) * $signed(input_fmap_92[7:0]) +
	( 11'sd 905) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18169) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10132) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12144) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6011) * $signed(input_fmap_97[7:0]) +
	( 11'sd 895) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11601) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14125) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8355) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11419) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18838) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2407) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8629) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4282) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12112) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12438) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18403) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17815) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13185) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17928) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4850) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29323) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8874) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24187) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 15'sd 15478) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1710) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6642) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31203) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27591) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29003) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16822) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28528) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23050) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6060) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25136) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1314) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32168) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20501) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_22[7:0]) +
	( 9'sd 176) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26021) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4715) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25668) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26943) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2192) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23878) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29959) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18219) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18291) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21072) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5210) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17755) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17603) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29033) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18113) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5625) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9056) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31187) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8211) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29212) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26337) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20234) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31673) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1896) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6572) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9428) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25140) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9261) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17095) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16060) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25674) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3409) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14900) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15117) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2927) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20148) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6809) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12730) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3698) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27947) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20352) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1070) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4684) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19808) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4841) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12534) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15478) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12422) * $signed(input_fmap_107[7:0]) +
	( 11'sd 951) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14898) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19134) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5875) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23778) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7553) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4743) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12637) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27605) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21931) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5087) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23828) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28016) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4222) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 16'sd 23390) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4415) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19530) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14230) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16982) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18044) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4975) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12157) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25248) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31728) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5710) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_21[7:0]) +
	( 9'sd 248) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1875) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28871) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31789) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24436) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11047) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24091) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11657) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4772) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28122) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_33[7:0]) +
	( 7'sd 58) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5725) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17050) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21279) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21272) * $signed(input_fmap_43[7:0]) +
	( 10'sd 350) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27830) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9827) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18824) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5390) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25427) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8224) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31283) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28506) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26855) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15181) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2754) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6857) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26701) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10502) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11219) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21912) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7398) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1129) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29209) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22690) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24628) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32689) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11609) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7645) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3634) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4346) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13434) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22433) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24761) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12464) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3860) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12015) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9688) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7646) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15527) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25722) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3838) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9799) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15819) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30375) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3490) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19983) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7767) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18873) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27483) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29548) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27844) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29932) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4136) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32111) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 15'sd 10662) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30415) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27313) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29454) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13928) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15987) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31996) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29270) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19580) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5985) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2363) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15834) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25743) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7891) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28041) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5407) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27082) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8886) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6709) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31011) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17766) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15632) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_37[7:0]) +
	( 11'sd 1006) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16833) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20556) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9363) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29022) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31572) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9003) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4599) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1363) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19351) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25314) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14980) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3113) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15131) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22120) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12365) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3029) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18752) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9216) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18005) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29564) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20245) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_85[7:0]) +
	( 10'sd 428) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7815) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31810) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14365) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11472) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6829) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20081) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10626) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14551) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6388) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13854) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24295) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21408) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16972) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8718) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31589) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10615) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7140) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28716) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28780) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6186) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4392) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2694) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10766) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29147) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10025) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17250) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22395) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31303) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24810) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 14'sd 4194) * $signed(input_fmap_0[7:0]) +
	( 10'sd 473) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30447) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_4[7:0]) +
	( 11'sd 976) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31394) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6593) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7512) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22347) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24504) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11725) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27857) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31056) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10994) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26514) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17981) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25031) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11640) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15364) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20925) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20573) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15203) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15864) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12142) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1070) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13061) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16049) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9478) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13862) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27610) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2051) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32362) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6969) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22665) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20215) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14433) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20149) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28860) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_67[7:0]) +
	( 10'sd 486) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14117) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5892) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8818) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11486) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5235) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12694) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28448) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7800) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16136) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11085) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22897) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31336) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8522) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22724) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18390) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4613) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17440) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27981) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27177) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7647) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10936) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26651) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23082) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_104[7:0]) +
	( 11'sd 761) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10779) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29196) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28158) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24506) * $signed(input_fmap_110[7:0]) +
	( 8'sd 71) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22080) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15567) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31542) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24407) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9922) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7665) * $signed(input_fmap_118[7:0]) +
	( 11'sd 964) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1154) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28997) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3950) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31769) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6429) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19524) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 14'sd 5686) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22310) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25329) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27454) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18347) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_8[7:0]) +
	( 11'sd 575) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25375) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2906) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28325) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6758) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22912) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23409) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6488) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25019) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31548) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2576) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24115) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_29[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24861) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10583) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20505) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14661) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10520) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29516) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2817) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11649) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28197) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29261) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7198) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29656) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9130) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25287) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19738) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23112) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3451) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32168) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32693) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1763) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10604) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31797) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15815) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25061) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30818) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23538) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21850) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18103) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15676) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17636) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21754) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27447) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24787) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12971) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18766) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5098) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6229) * $signed(input_fmap_85[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2972) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20508) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12164) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13854) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16914) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21549) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27324) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3768) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12218) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32445) * $signed(input_fmap_103[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11785) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31155) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19682) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23861) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26694) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24784) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23090) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9045) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14495) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26842) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23708) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22608) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24308) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17232) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_124[7:0]) +
	( 9'sd 214) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1169) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 15'sd 15801) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24185) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7608) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9186) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3578) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12037) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13358) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5807) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4534) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22493) * $signed(input_fmap_14[7:0]) +
	( 10'sd 380) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18457) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21518) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4932) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18227) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8182) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31793) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_28[7:0]) +
	( 12'sd 2032) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13865) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9863) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4098) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1432) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5543) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28672) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13100) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29482) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16390) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13034) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28987) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24384) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22023) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3891) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20887) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24844) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11241) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13195) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_57[7:0]) +
	( 14'sd 8028) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16790) * $signed(input_fmap_60[7:0]) +
	( 11'sd 587) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2144) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8706) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31520) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32072) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30051) * $signed(input_fmap_68[7:0]) +
	( 8'sd 83) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24283) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27837) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16805) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26183) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10177) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17736) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5659) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24288) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18399) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20933) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3946) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12191) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22844) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3874) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21911) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3425) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17479) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5964) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30950) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6402) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24505) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12797) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21632) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11086) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10991) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18714) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18540) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10967) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2996) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12372) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24857) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29777) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27648) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10436) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26063) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 16'sd 29532) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12618) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_2[7:0]) +
	( 10'sd 288) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7302) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29343) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12716) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20137) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9323) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25045) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24329) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11478) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_14[7:0]) +
	( 10'sd 303) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17975) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5860) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17479) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16058) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23352) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16122) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13124) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5181) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13827) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24367) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5472) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10053) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32251) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15207) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3858) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19236) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22446) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6410) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18884) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20576) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2052) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28966) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13510) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2522) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1863) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6979) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29796) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28942) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28824) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16148) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17804) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31497) * $signed(input_fmap_65[7:0]) +
	( 7'sd 46) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7380) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14172) * $signed(input_fmap_68[7:0]) +
	( 15'sd 16354) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5293) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24566) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21148) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19577) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6081) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21942) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18576) * $signed(input_fmap_78[7:0]) +
	( 11'sd 835) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9587) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18552) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29459) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32335) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17063) * $signed(input_fmap_84[7:0]) +
	( 11'sd 995) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6271) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9065) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26136) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13919) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21416) * $signed(input_fmap_93[7:0]) +
	( 9'sd 224) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5598) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9524) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1827) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14711) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31230) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11661) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3942) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27963) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11991) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19792) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18447) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32623) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25643) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29584) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_120[7:0]) +
	( 10'sd 477) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28057) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8217) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16542) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13048) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13733) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3174) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 16'sd 28203) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13719) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19937) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22355) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15285) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_7[7:0]) +
	( 10'sd 424) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4709) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23189) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5164) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31666) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7343) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22529) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14113) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6205) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20731) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15356) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11483) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16219) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10077) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29906) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23861) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10755) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18979) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10422) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13044) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11508) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18498) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5194) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21188) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22967) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32366) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1283) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31020) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18863) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22711) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9697) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17953) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26033) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14302) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9642) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16642) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2924) * $signed(input_fmap_78[7:0]) +
	( 11'sd 958) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25202) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26018) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14154) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17701) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11640) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7614) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23046) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26327) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31478) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6003) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14352) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17201) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2895) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27300) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16243) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15467) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16936) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6716) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18247) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20583) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13554) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1570) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23401) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18204) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29173) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5775) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26384) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19065) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21101) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4569) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2820) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_122[7:0]) +
	( 10'sd 434) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5756) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1427) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26883) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 11'sd 527) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14573) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16125) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25114) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24504) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15407) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16965) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12569) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31601) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25388) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26817) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21354) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17540) * $signed(input_fmap_22[7:0]) +
	( 10'sd 389) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23276) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26134) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1306) * $signed(input_fmap_29[7:0]) +
	( 13'sd 4046) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14896) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19257) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16163) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18277) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23112) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29944) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20975) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6011) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30786) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18129) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11035) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25304) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2304) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3400) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21359) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25990) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32374) * $signed(input_fmap_48[7:0]) +
	( 11'sd 679) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24856) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3128) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22727) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20053) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24548) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29810) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4917) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29476) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25959) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18394) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7997) * $signed(input_fmap_65[7:0]) +
	( 11'sd 779) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6254) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_68[7:0]) +
	( 15'sd 16336) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17988) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19853) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21093) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22713) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22763) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23442) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14528) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27135) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19163) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9251) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19860) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15117) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9520) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2598) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1287) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13901) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12803) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3455) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20962) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24920) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23598) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19879) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8235) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26422) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30054) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22609) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11207) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32282) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3129) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3518) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10517) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2199) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2809) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24923) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16669) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18738) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31913) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21167) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18585) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32392) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26042) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5866) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30937) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23714) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 14'sd 4421) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_1[7:0]) +
	( 11'sd 931) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6483) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6888) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4674) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22677) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31663) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1625) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12873) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16160) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27469) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31148) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15595) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16231) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2285) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26440) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6028) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5980) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26805) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31763) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19099) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7347) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25580) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4477) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18465) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29309) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23828) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30256) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23179) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29918) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1910) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13057) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18821) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26490) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_54[7:0]) +
	( 7'sd 57) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26190) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5546) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7284) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27570) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20205) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19779) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32085) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30838) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30690) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3134) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26203) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15775) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12724) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6264) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29554) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32655) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12783) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7258) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16871) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12114) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2208) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31919) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11169) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8342) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26305) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7610) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19794) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6350) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23225) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30151) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7832) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30526) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6818) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7371) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22803) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14013) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8745) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26779) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24053) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27518) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20539) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15204) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13115) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12518) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30260) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28992) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20879) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3917) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2233) * $signed(input_fmap_122[7:0]) +
	( 6'sd 30) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2208) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26907) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 14'sd 4921) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8268) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22147) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17892) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26470) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1894) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11776) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26246) * $signed(input_fmap_8[7:0]) +
	( 12'sd 2017) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13976) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2956) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4670) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1585) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11060) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16275) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24871) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14359) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16136) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4724) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32353) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14459) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26042) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17663) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1121) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18961) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4926) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13077) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8581) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7681) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31706) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17071) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6881) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25465) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_52[7:0]) +
	( 11'sd 943) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29213) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16395) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29678) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26408) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23135) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6812) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12243) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26907) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6586) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22936) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5528) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30546) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25127) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1583) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7259) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17897) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9623) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10245) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12267) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8979) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16211) * $signed(input_fmap_88[7:0]) +
	( 11'sd 961) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12578) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9620) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12540) * $signed(input_fmap_92[7:0]) +
	( 11'sd 519) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32305) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21932) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26188) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22146) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29276) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13056) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28681) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29088) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32662) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4354) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18483) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11215) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16700) * $signed(input_fmap_116[7:0]) +
	( 11'sd 615) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29731) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19136) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1607) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26638) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15380) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 16'sd 21044) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2948) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13788) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28517) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21330) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32031) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19519) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28008) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23429) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31194) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13744) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31891) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24583) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24383) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24646) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5469) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5492) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18429) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_22[7:0]) +
	( 11'sd 574) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5350) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24324) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19629) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11004) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13457) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21141) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16360) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25269) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4423) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1317) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26974) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16143) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1166) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4964) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2919) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_48[7:0]) +
	( 10'sd 417) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24307) * $signed(input_fmap_51[7:0]) +
	( 5'sd 15) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10009) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19427) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3359) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11788) * $signed(input_fmap_57[7:0]) +
	( 9'sd 252) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31162) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14997) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15741) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14022) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31137) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4272) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1709) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18138) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6365) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30869) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13022) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5902) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31208) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1903) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22053) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1461) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29741) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25795) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18169) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_92[7:0]) +
	( 11'sd 937) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11854) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27529) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20321) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6721) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9206) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10953) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21471) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14193) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5859) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27854) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1176) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15519) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27360) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20250) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13668) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_113[7:0]) +
	( 13'sd 4067) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10177) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13646) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10227) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25873) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28032) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29408) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 16'sd 27680) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17870) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8727) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15054) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10171) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16271) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17723) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1543) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16226) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29680) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17512) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13463) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22279) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2532) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2578) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1031) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32587) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5869) * $signed(input_fmap_28[7:0]) +
	( 11'sd 912) * $signed(input_fmap_29[7:0]) +
	( 10'sd 417) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25826) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1823) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6773) * $signed(input_fmap_34[7:0]) +
	( 11'sd 847) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20216) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21969) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10433) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8864) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8856) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22362) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15409) * $signed(input_fmap_45[7:0]) +
	( 14'sd 8032) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15447) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20621) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17965) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11877) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17808) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12829) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7669) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10099) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21909) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23339) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6750) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13821) * $signed(input_fmap_70[7:0]) +
	( 10'sd 413) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15828) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31675) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19234) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26403) * $signed(input_fmap_79[7:0]) +
	( 10'sd 358) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2077) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23644) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5741) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23253) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7983) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27171) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32588) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12023) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31808) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3504) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14973) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5849) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13067) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29663) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1206) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_110[7:0]) +
	( 11'sd 889) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13668) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21244) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2514) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_124[7:0]) +
	( 11'sd 584) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25821) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 9'sd 202) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31324) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27003) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14186) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27291) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25580) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8745) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9501) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13921) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19290) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25188) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21277) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7567) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19345) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11158) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10265) * $signed(input_fmap_27[7:0]) +
	( 10'sd 466) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30487) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19248) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14309) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21521) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19306) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15153) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30787) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3691) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14393) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10649) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3790) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1100) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18003) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16143) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24177) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2398) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18979) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30197) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20194) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30002) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27042) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2822) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29381) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29688) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31308) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3389) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12713) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24645) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27570) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30493) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5125) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3386) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24134) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2699) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26943) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30450) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4829) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15683) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11306) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3974) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29859) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8381) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21242) * $signed(input_fmap_99[7:0]) +
	( 7'sd 42) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7415) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8882) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3169) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28202) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16313) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27530) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5079) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17379) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15646) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18643) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32217) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2126) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13771) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 13'sd 2302) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17126) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16607) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13778) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4949) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_5[7:0]) +
	( 11'sd 844) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4222) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25594) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16889) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2100) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21400) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25283) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6854) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7027) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27849) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20187) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19386) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3555) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3236) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16970) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18602) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10020) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20521) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1483) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31305) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9418) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13068) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20386) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29574) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17829) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13479) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16480) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14912) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27747) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3437) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12033) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17018) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30294) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23523) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11415) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11625) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4427) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_67[7:0]) +
	( 11'sd 999) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10217) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29935) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20800) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8829) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5489) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29367) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21615) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24824) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18044) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5202) * $signed(input_fmap_84[7:0]) +
	( 11'sd 1010) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8236) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28587) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10581) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27287) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7456) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14698) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3398) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25398) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6515) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26559) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13417) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21713) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1498) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16601) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29800) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14452) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6495) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24536) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27584) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14893) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23587) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11095) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4485) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27031) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22382) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23102) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 16'sd 24528) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5041) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18170) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31619) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28123) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25131) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26723) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1345) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31023) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23217) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22430) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5595) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17653) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25711) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27648) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31635) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30640) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6385) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28865) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7691) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14644) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32339) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1328) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25329) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13192) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21970) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25377) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8213) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6224) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24326) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11876) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2255) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21374) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15664) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6327) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4315) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31772) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6560) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7160) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30682) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31313) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20576) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30764) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15037) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13487) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20998) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12117) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24154) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11047) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17066) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25323) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31357) * $signed(input_fmap_86[7:0]) +
	( 9'sd 210) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9999) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17149) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6721) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20858) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_96[7:0]) +
	( 9'sd 255) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5341) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28311) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5811) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12299) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9876) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5057) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1978) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20623) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6622) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30433) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25114) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12995) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29031) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22489) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18565) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10498) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5765) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22722) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 12'sd 1048) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3480) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31592) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19335) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29403) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1437) * $signed(input_fmap_6[7:0]) +
	( 11'sd 736) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31790) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10484) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12943) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23601) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31991) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4525) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10506) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20377) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13164) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9703) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13344) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13544) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23787) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18920) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1264) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1942) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14735) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24699) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32332) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16428) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15874) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10140) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11368) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2546) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2537) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26705) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_55[7:0]) +
	( 11'sd 649) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17076) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26777) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3104) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15355) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16745) * $signed(input_fmap_64[7:0]) +
	( 11'sd 767) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12594) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4570) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11948) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10704) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17044) * $signed(input_fmap_72[7:0]) +
	( 10'sd 468) * $signed(input_fmap_73[7:0]) +
	( 11'sd 793) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31557) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11103) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3333) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23702) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8979) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24274) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13376) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28504) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1401) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7796) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20217) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28998) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20854) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31055) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2715) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21160) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21628) * $signed(input_fmap_101[7:0]) +
	( 10'sd 450) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6589) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17458) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29209) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15957) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11478) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9055) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13955) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10273) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11173) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8100) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22713) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3860) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26484) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3473) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12705) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12263) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14218) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 27093) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11084) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24722) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9427) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11753) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14913) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4870) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32299) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26642) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6330) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25757) * $signed(input_fmap_18[7:0]) +
	( 11'sd 633) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30098) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19927) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7851) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6103) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9915) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19392) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2712) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7320) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22380) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19349) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18340) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31376) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1645) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20742) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12396) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17152) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_46[7:0]) +
	( 11'sd 849) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25496) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28189) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25951) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14792) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26347) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6495) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31024) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5919) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1542) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18045) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19937) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21914) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14883) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6331) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_74[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1926) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27350) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31361) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21892) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21548) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27638) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26145) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23107) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29302) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10145) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31674) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11913) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3844) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31716) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9749) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22199) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24429) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2331) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29563) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16640) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21969) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29862) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9376) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31083) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12767) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25303) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24692) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26860) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2376) * $signed(input_fmap_126[7:0]) +
	( 6'sd 17) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 16'sd 28441) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16127) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1623) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27872) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_5[7:0]) +
	( 11'sd 961) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24790) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19659) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15388) * $signed(input_fmap_9[7:0]) +
	( 10'sd 444) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14034) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3199) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1997) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9013) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1152) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14582) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32163) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2289) * $signed(input_fmap_25[7:0]) +
	( 9'sd 174) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27596) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7686) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5643) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29087) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16105) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31231) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15403) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5089) * $signed(input_fmap_39[7:0]) +
	( 11'sd 998) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1691) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30308) * $signed(input_fmap_42[7:0]) +
	( 11'sd 755) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25429) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12653) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13920) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2096) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9063) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1831) * $signed(input_fmap_54[7:0]) +
	( 11'sd 691) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12245) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5572) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8228) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18753) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29791) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23752) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4552) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4392) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13336) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21978) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14809) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15855) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3433) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23126) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8466) * $signed(input_fmap_80[7:0]) +
	( 9'sd 159) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3135) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7144) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29387) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1325) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25306) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18877) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12208) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11251) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19736) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21504) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21501) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14792) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10710) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15376) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28915) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13907) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8982) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12444) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_101[7:0]) +
	( 6'sd 26) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21505) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19219) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25513) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17982) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15906) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21513) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30085) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6124) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10282) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1349) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31884) * $signed(input_fmap_115[7:0]) +
	( 11'sd 696) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11731) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28128) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26565) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27920) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29688) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16868) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19009) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 16'sd 28985) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4932) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28458) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11248) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5716) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32735) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15958) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1128) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22362) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2423) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4412) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16330) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17083) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3910) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27573) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14334) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18378) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29417) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32204) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2533) * $signed(input_fmap_25[7:0]) +
	( 11'sd 828) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14044) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23217) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25719) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6390) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32706) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22219) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8359) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13408) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14347) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29640) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8605) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10962) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4218) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30595) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16433) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26754) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29407) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26302) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17302) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29003) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22282) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23948) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24441) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5787) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26302) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26415) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21365) * $signed(input_fmap_72[7:0]) +
	( 10'sd 491) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5647) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17062) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23677) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21298) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5061) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15750) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28391) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_86[7:0]) +
	( 10'sd 281) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3106) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13490) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22668) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16631) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24531) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9163) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29979) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7804) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10803) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11549) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17552) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12757) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32182) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20748) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22983) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3341) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14181) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26516) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5033) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15583) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17636) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29683) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23165) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4878) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25832) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2730) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3180) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31390) * $signed(input_fmap_121[7:0]) +
	( 9'sd 171) * $signed(input_fmap_122[7:0]) +
	( 13'sd 4066) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3298) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7031) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26308) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 14'sd 6352) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5140) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19181) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4297) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26312) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29741) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12970) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12594) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11742) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30121) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21125) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27337) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18954) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5316) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26783) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20878) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23109) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27209) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21323) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19392) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7482) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10116) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3061) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29284) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5914) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26771) * $signed(input_fmap_38[7:0]) +
	( 11'sd 637) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26098) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22366) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5083) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18372) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32628) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7422) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22028) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20032) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11733) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7737) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24494) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24087) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15799) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15320) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19647) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19183) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13065) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20918) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28992) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22942) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20298) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16786) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30071) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31576) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12889) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14209) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22242) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22684) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12647) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26227) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27326) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28234) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29236) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23423) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27423) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9068) * $signed(input_fmap_87[7:0]) +
	( 10'sd 435) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30640) * $signed(input_fmap_91[7:0]) +
	( 12'sd 2034) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29090) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3439) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5521) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4362) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29030) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13903) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21195) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29134) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16011) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7212) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32007) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_113[7:0]) +
	( 11'sd 595) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2195) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28338) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2223) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5926) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1084) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31366) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19312) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1865) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26538) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9286) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 16'sd 17136) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11522) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21149) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23258) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24288) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24275) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20743) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11417) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22321) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1221) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30239) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22751) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32352) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14172) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7807) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20666) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10591) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1318) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24230) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16566) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24892) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18206) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25823) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10747) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19151) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31628) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26892) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4166) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6433) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26262) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26214) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22653) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10654) * $signed(input_fmap_49[7:0]) +
	( 11'sd 922) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20277) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4226) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20833) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28560) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28752) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2954) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7170) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31190) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_62[7:0]) +
	( 10'sd 300) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10588) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30507) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30167) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14999) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32552) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6272) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25143) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27121) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25030) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18888) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4317) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29920) * $signed(input_fmap_89[7:0]) +
	( 7'sd 50) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7018) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25071) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25864) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1786) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5965) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1836) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8687) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23911) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14133) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1076) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24767) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28752) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11234) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27149) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12356) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17867) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5220) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10928) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10917) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13108) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18868) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25895) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1176) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24448) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4500) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23957) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30261) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32346) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23914) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12167) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29578) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22091) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 15'sd 15604) * $signed(input_fmap_0[7:0]) +
	( 6'sd 27) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22419) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29139) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25678) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3342) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24977) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8858) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24066) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21464) * $signed(input_fmap_13[7:0]) +
	( 11'sd 899) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12585) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22426) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15099) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22407) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30555) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26862) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6199) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27030) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17896) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11765) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14746) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13938) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1463) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22521) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19199) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1506) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30972) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11999) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8337) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_45[7:0]) +
	( 10'sd 443) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28455) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6528) * $signed(input_fmap_48[7:0]) +
	( 10'sd 459) * $signed(input_fmap_49[7:0]) +
	( 10'sd 342) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18832) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3378) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26565) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12664) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1609) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18474) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30484) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4494) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20983) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10374) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13812) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9468) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29538) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17650) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17562) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9914) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1784) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25435) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10559) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4505) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25328) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_84[7:0]) +
	( 8'sd 66) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7928) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29427) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16566) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23299) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12490) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20092) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9686) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_100[7:0]) +
	( 10'sd 359) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32521) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20156) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15649) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3125) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8556) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18557) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3610) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29662) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4545) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22294) * $signed(input_fmap_115[7:0]) +
	( 9'sd 206) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17079) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28054) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11834) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15224) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24330) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 16'sd 29894) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16022) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21354) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20443) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25624) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4719) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9920) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27421) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9108) * $signed(input_fmap_14[7:0]) +
	( 7'sd 59) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13418) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26234) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12683) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26731) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22860) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9559) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13635) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15225) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32245) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19522) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3062) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19616) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29276) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28478) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2936) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8626) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21467) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1661) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10067) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7383) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7518) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5474) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16568) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23819) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15894) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19904) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_72[7:0]) +
	( 9'sd 157) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30478) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25504) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28776) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_81[7:0]) +
	( 10'sd 313) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8848) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2452) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8498) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3173) * $signed(input_fmap_87[7:0]) +
	( 11'sd 795) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22863) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23447) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31875) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26045) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32318) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2804) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17109) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_98[7:0]) +
	( 11'sd 891) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25328) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30452) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28643) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7200) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4523) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9675) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19783) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27791) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14811) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23331) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11607) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6258) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10683) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3601) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26168) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 16'sd 31022) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12553) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26672) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6794) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12787) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8912) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29469) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13374) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_10[7:0]) +
	( 13'sd 4082) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9658) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32303) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18775) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10988) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30415) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9842) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22240) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22059) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11324) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31536) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10396) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15244) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32200) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24194) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2543) * $signed(input_fmap_34[7:0]) +
	( 11'sd 598) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4909) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13044) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23880) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7182) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7191) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20205) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10243) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11712) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16213) * $signed(input_fmap_52[7:0]) +
	( 11'sd 699) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30825) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14770) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3747) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_60[7:0]) +
	( 12'sd 2030) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30462) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15342) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28581) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26344) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7758) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12890) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13621) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9307) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_73[7:0]) +
	( 11'sd 965) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28213) * $signed(input_fmap_76[7:0]) +
	( 13'sd 4048) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15930) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13216) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16584) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26297) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7054) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8260) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9585) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7661) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3500) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13546) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15446) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3251) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24962) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18640) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12732) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30947) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26593) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28083) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17993) * $signed(input_fmap_100[7:0]) +
	( 7'sd 61) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3873) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5571) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31889) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7626) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22419) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7126) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12027) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20355) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32588) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30215) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19547) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24603) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14422) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 16'sd 21952) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11510) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1951) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7229) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24384) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29852) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11290) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27132) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18980) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4950) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18729) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26452) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18048) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31464) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19380) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23717) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6855) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6043) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20618) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20746) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27200) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22639) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_29[7:0]) +
	( 11'sd 591) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16092) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12096) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11128) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31629) * $signed(input_fmap_36[7:0]) +
	( 11'sd 992) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15276) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12968) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8350) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16436) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21260) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23781) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30522) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8687) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5162) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32041) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1402) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30092) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23986) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32326) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9615) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22870) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31805) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29245) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3343) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6693) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23934) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8161) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12239) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27020) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25519) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_71[7:0]) +
	( 11'sd 932) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20014) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26643) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17991) * $signed(input_fmap_75[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31278) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18897) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31024) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12745) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4200) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30859) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_85[7:0]) +
	( 6'sd 29) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28211) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30607) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14074) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12602) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26418) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6641) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12174) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15092) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27097) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29634) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29745) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13918) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9074) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24557) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6635) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1028) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_112[7:0]) +
	( 9'sd 130) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28832) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2088) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13821) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21554) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8540) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21304) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 12'sd 1272) * $signed(input_fmap_0[7:0]) +
	( 11'sd 768) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18225) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12530) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11059) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10410) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16584) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4933) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23184) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22719) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27245) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26964) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12175) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28079) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15806) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31183) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21358) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32236) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9008) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16405) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10754) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25905) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5427) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25713) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20739) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31910) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19860) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11362) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13752) * $signed(input_fmap_45[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_47[7:0]) +
	( 10'sd 472) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6460) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10501) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8048) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1048) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30514) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24534) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8827) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10464) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4535) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15398) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5119) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14218) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31300) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23890) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20574) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4765) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31748) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23124) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15189) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10436) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26753) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26739) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15375) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23969) * $signed(input_fmap_80[7:0]) +
	( 8'sd 111) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9616) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_85[7:0]) +
	( 11'sd 980) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27962) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6266) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14458) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20157) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5486) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2142) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16233) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29617) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20901) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19536) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9423) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31827) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23970) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26993) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1604) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22780) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_108[7:0]) +
	( 9'sd 252) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17087) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8452) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27907) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9091) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21929) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9103) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6437) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_122[7:0]) +
	( 9'sd 210) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2170) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7157) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26028) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 11'sd 596) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13145) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26770) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28298) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7636) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20761) * $signed(input_fmap_16[7:0]) +
	( 11'sd 804) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28833) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14948) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24661) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25370) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28078) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2660) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22534) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15792) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26609) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16512) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15218) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18392) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_36[7:0]) +
	( 11'sd 606) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21701) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20262) * $signed(input_fmap_40[7:0]) +
	( 11'sd 550) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32052) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27897) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9544) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24137) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27345) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19113) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27931) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27732) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31450) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24949) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27161) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22695) * $signed(input_fmap_62[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29546) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17338) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7729) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12163) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26130) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10904) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29783) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9896) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27259) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31057) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15650) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3152) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26413) * $signed(input_fmap_86[7:0]) +
	( 8'sd 116) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11804) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24305) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27276) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32540) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5929) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31090) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30628) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32293) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16419) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2656) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25262) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7997) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8298) * $signed(input_fmap_111[7:0]) +
	( 11'sd 750) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17847) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6241) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7873) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17656) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31207) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2384) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12657) * $signed(input_fmap_122[7:0]) +
	( 11'sd 616) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12919) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16599) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20111) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 16'sd 25069) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29558) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2670) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4113) * $signed(input_fmap_3[7:0]) +
	( 9'sd 220) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27031) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25621) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5864) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26653) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30997) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28915) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3854) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8959) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7457) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17466) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5737) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32727) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8606) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4476) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15611) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6557) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23678) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30581) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26560) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8894) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28185) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22862) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18048) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6054) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3477) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3542) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18483) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18537) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28379) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1450) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15371) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24607) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_51[7:0]) +
	( 10'sd 419) * $signed(input_fmap_52[7:0]) +
	( 13'sd 4013) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8100) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18194) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19547) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12406) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26341) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1412) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32159) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16726) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17554) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25871) * $signed(input_fmap_71[7:0]) +
	( 10'sd 324) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16125) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17087) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1060) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23969) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14329) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1214) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5517) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2413) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31925) * $signed(input_fmap_88[7:0]) +
	( 7'sd 53) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25632) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11112) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30879) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8638) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16813) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1687) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5132) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1825) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25670) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14265) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9391) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26409) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10561) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32025) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10864) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18954) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21276) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32481) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26262) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3437) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14206) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19978) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22004) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16210) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23387) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3489) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 16'sd 22891) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19791) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5014) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14674) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24202) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15795) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32491) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9203) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10446) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3512) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13618) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30495) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22247) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9814) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17829) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3543) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27011) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16798) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19129) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28915) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12973) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3265) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8313) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22538) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28508) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10754) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21982) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21802) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31158) * $signed(input_fmap_40[7:0]) +
	( 11'sd 792) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24524) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9401) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3300) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3665) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_50[7:0]) +
	( 9'sd 153) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24623) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7386) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4853) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21459) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15889) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6625) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4299) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4923) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9357) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21259) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17879) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17267) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27033) * $signed(input_fmap_74[7:0]) +
	( 11'sd 985) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22035) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11825) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29295) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15386) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23763) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13302) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18067) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28330) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8972) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19756) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4708) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3129) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20541) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11231) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31896) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21505) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20558) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12386) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6581) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13098) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3515) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13160) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27920) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1390) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28759) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4143) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11713) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30752) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9941) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29553) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9129) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20323) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32754) * $signed(input_fmap_124[7:0]) +
	( 8'sd 99) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20526) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 16'sd 19537) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23179) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29749) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6311) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26472) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19977) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15724) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31423) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12964) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25761) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19222) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30605) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8063) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31235) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30477) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10794) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5893) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26098) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32765) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6087) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19427) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23476) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16322) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15046) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6237) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25250) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26546) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16710) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10224) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30834) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27200) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3722) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19013) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30358) * $signed(input_fmap_43[7:0]) +
	( 13'sd 4083) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17807) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24119) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31608) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26762) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11167) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17366) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16269) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31404) * $signed(input_fmap_61[7:0]) +
	( 7'sd 46) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2751) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3834) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7045) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29063) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1679) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6798) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10982) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13522) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4431) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8817) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14528) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27297) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7358) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8570) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24729) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18258) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24757) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13977) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16210) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20968) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4120) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17396) * $signed(input_fmap_92[7:0]) +
	( 9'sd 205) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32291) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10336) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17272) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14862) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10306) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20083) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22769) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20639) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7263) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20126) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29219) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26835) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27770) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18891) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32572) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_124[7:0]) +
	( 9'sd 240) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3682) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 16'sd 17368) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16749) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5141) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28505) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21782) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10307) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19319) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27401) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2917) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12609) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29673) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8600) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_22[7:0]) +
	( 8'sd 110) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10659) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13619) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24119) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25143) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28956) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19121) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3785) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21027) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24708) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28149) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16377) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22916) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32557) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19747) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21810) * $signed(input_fmap_44[7:0]) +
	( 14'sd 8171) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1990) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17486) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_48[7:0]) +
	( 11'sd 919) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26989) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23990) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12260) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16146) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17655) * $signed(input_fmap_55[7:0]) +
	( 8'sd 83) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15690) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20432) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1127) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22936) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7214) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13271) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26838) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24221) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24100) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20819) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23432) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24030) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17241) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3110) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4567) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3439) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22936) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29945) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7283) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28382) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13663) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13525) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14586) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14603) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6440) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3229) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19980) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1856) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20648) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6972) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21329) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18078) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18687) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5879) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10044) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8973) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24639) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32643) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22536) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3343) * $signed(input_fmap_111[7:0]) +
	( 14'sd 8076) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25692) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31776) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11265) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5626) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29411) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23951) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24680) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15814) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 13'sd 3089) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14753) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12252) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20242) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17900) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18979) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7832) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16986) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12398) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4778) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7475) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10621) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7229) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29081) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3412) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27811) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7388) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11999) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22530) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7956) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31463) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14023) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12651) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13536) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26972) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25576) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20787) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22322) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24785) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30362) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12868) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5563) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23722) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25615) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30122) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18042) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18955) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24329) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4554) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2792) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_54[7:0]) +
	( 7'sd 38) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30116) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29252) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13900) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30253) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4597) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28002) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16206) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18610) * $signed(input_fmap_65[7:0]) +
	( 10'sd 386) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10126) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27556) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13944) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27590) * $signed(input_fmap_74[7:0]) +
	( 14'sd 8055) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25732) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29222) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6142) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9648) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32441) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1898) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5693) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9113) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29552) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32005) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4954) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1407) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16450) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24074) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19655) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30288) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22298) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20879) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16167) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6536) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22973) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_113[7:0]) +
	( 11'sd 782) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3246) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18524) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14383) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32175) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14816) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27386) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8425) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13313) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5272) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25203) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 16'sd 29620) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23957) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19253) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16099) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1693) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20628) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2433) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19282) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17576) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17027) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10345) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27712) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15343) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27449) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27731) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20595) * $signed(input_fmap_21[7:0]) +
	( 9'sd 212) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17112) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12056) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2934) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7768) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8298) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6331) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1398) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7758) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25654) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6668) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17974) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27646) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21784) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22861) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8387) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12827) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1381) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10485) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16574) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13933) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15224) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11402) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1726) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25158) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22313) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_58[7:0]) +
	( 9'sd 193) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10240) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1447) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15222) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8930) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4299) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8349) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19418) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17213) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28922) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13288) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5267) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18237) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19488) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21489) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15400) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5569) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21290) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31067) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15273) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7687) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26506) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5931) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27751) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11728) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31576) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18373) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12960) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29655) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17872) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13448) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7673) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3099) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5501) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20230) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21485) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26451) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18182) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2661) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12921) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31877) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30663) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16660) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21923) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32209) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9553) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8453) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18618) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 16'sd 18457) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4252) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4428) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7334) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7686) * $signed(input_fmap_4[7:0]) +
	( 9'sd 224) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3488) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22529) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17738) * $signed(input_fmap_10[7:0]) +
	( 10'sd 462) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17725) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1173) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9650) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30783) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8960) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_21[7:0]) +
	( 14'sd 8090) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25010) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26010) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8906) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25489) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22560) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13824) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30656) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18653) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7768) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24533) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_37[7:0]) +
	( 9'sd 145) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9657) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25871) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10837) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20113) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13653) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25990) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26874) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1527) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6651) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32338) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21849) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24160) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13789) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5199) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19749) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17215) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9312) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32164) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14261) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7460) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19286) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16003) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9102) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29395) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1229) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19525) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14739) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12815) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31568) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27092) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27733) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14363) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10649) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4200) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3699) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9684) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25704) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9949) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10915) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13149) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27638) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1431) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12000) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19427) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21434) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16589) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30686) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4331) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20516) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16271) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1255) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12269) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27592) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30242) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12024) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15993) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23529) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30747) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 10'sd 431) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19951) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4474) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20012) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15800) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9501) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29228) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32079) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5246) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22045) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8594) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13376) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28502) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18745) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11786) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8729) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4206) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1798) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10701) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12517) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22262) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17799) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8008) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1885) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19673) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4650) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20035) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26323) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3385) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20136) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11642) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11292) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3725) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13445) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12931) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15301) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12560) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21090) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14339) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6528) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21420) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6049) * $signed(input_fmap_60[7:0]) +
	( 11'sd 936) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20042) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27901) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27683) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32105) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14725) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31063) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23623) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21302) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1363) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24757) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22804) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16936) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28341) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8369) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21850) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2898) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15089) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28072) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11578) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19109) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8474) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16150) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3430) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18316) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5783) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14563) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21264) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20555) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10187) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1567) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9363) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25586) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11763) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14766) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3124) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_122[7:0]) +
	( 8'sd 107) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26000) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4999) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28655) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 14'sd 4893) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31511) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16857) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13502) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25851) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19342) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21304) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14393) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23190) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25098) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10699) * $signed(input_fmap_15[7:0]) +
	( 11'sd 760) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32285) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11842) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18773) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10530) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5717) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32102) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7299) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28534) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_30[7:0]) +
	( 14'sd 8156) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9512) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20251) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5536) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25581) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22025) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4827) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28756) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16605) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25208) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4644) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_48[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9209) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23426) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21841) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13709) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31132) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8221) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13751) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14378) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9367) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17949) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30746) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22509) * $signed(input_fmap_69[7:0]) +
	( 10'sd 435) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24315) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2973) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21520) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7110) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20541) * $signed(input_fmap_80[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29386) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7662) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28813) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_91[7:0]) +
	( 11'sd 952) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10760) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4465) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17240) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22695) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14632) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15809) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6340) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21916) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26536) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10672) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16542) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26672) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19634) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31685) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15637) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10582) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28314) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14906) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11697) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26001) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8693) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9199) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 16'sd 29741) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19493) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6481) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10520) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2598) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8563) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14624) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29891) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17567) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10462) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9263) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9077) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5789) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17258) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30870) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29684) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15971) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30520) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9906) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5980) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8692) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3708) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9994) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31990) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22944) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8586) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27151) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32287) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5539) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22509) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28901) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8417) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17795) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9707) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5339) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7670) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5706) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15103) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17933) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27698) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6216) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21484) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15483) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27317) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3831) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27732) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19366) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28390) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3049) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8818) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19276) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19202) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11949) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23245) * $signed(input_fmap_86[7:0]) +
	( 11'sd 976) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32456) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20291) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13438) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9641) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27006) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7758) * $signed(input_fmap_95[7:0]) +
	( 11'sd 808) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21720) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22265) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24951) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32236) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24746) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31543) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21358) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30314) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7237) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27630) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1317) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19612) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12465) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29300) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7936) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13237) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4464) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 15'sd 14406) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32705) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17963) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25316) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4297) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2126) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10216) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9495) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23164) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25634) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4182) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23871) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6518) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29625) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27115) * $signed(input_fmap_26[7:0]) +
	( 11'sd 576) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29906) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14113) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1524) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9180) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27880) * $signed(input_fmap_35[7:0]) +
	( 11'sd 553) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15295) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10258) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22334) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_40[7:0]) +
	( 9'sd 224) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19774) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16155) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_44[7:0]) +
	( 13'sd 4016) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11655) * $signed(input_fmap_49[7:0]) +
	( 10'sd 302) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28441) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7995) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3172) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3635) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3069) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20242) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28756) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29975) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13789) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20295) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2863) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11352) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31730) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23474) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10987) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31608) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7480) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4759) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6970) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28905) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24845) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17323) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9675) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30014) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31137) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10761) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29965) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17338) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14812) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_102[7:0]) +
	( 12'sd 2026) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14853) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5837) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27944) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6001) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1985) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15208) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6763) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21708) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16989) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28485) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31222) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30145) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21729) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2255) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28341) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 15'sd 8981) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16569) * $signed(input_fmap_1[7:0]) +
	( 10'sd 492) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28151) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9712) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15972) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17296) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1232) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25073) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11759) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29536) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28128) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30713) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8529) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23026) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31448) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9232) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21207) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25184) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25091) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17608) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9905) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29791) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21929) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4179) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8660) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30284) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29834) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14311) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18947) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21621) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3134) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30428) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_50[7:0]) +
	( 9'sd 171) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30935) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9041) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28780) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13512) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12676) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31231) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2278) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31409) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17434) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15492) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16910) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28386) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19813) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13536) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22594) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24139) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_86[7:0]) +
	( 11'sd 782) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14793) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9800) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17645) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8724) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21477) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13192) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9730) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19434) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27827) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4250) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9840) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13776) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16805) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23996) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3366) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24619) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10463) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11541) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24120) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18085) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 16'sd 25468) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30875) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12158) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17741) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18875) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12369) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21551) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8343) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12102) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15505) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13658) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21253) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16751) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5128) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8469) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24286) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20773) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18171) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26482) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31951) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7453) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12252) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25169) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14847) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20638) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21352) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10912) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18767) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15156) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8400) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5524) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2433) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18030) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6421) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25960) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21867) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10938) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9105) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26452) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14055) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9137) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11156) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5896) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29490) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12510) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4223) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28488) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6816) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8588) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24034) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9071) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27849) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7303) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4731) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31119) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18221) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8992) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29871) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32510) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26320) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18027) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24670) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14074) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13729) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9622) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17219) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5116) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20967) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13815) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30792) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28232) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24371) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12125) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14576) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7086) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18617) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6032) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30450) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6778) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32247) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19034) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 12'sd 1194) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20881) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15224) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19317) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19894) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1401) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19426) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19983) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25324) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20610) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23758) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7631) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22318) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11434) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26242) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32543) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25396) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8417) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4609) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21127) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20715) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31070) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27153) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19986) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7255) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2856) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8366) * $signed(input_fmap_38[7:0]) +
	( 11'sd 747) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27646) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4346) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5535) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5463) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3674) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32490) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15978) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12808) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22775) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25034) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22012) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2143) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_60[7:0]) +
	( 11'sd 611) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7444) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21348) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26083) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1641) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20236) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31754) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7308) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16782) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20209) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20656) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21918) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4378) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10442) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17213) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1900) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7662) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16100) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8045) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12747) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8897) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8882) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19452) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2236) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26929) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21154) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22227) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20609) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30527) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25818) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12234) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5395) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17328) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15117) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10078) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30472) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23835) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4972) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28572) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15937) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13628) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1558) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 14'sd 5799) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25545) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8376) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14409) * $signed(input_fmap_3[7:0]) +
	( 9'sd 197) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32549) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20080) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5198) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11758) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25354) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13319) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19294) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3945) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23141) * $signed(input_fmap_14[7:0]) +
	( 8'sd 106) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23703) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31732) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19537) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19402) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12313) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25258) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23447) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11958) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30942) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1287) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31890) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17354) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31416) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6057) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31056) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30987) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7529) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25444) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9134) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26474) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31710) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26723) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16080) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12917) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20506) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17238) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17971) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14899) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11541) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_52[7:0]) +
	( 9'sd 130) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31988) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13178) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25759) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24855) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14333) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21478) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12167) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30922) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20977) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15764) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4606) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25450) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17098) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15068) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32655) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28128) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10492) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13909) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20240) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10794) * $signed(input_fmap_85[7:0]) +
	( 8'sd 74) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21295) * $signed(input_fmap_88[7:0]) +
	( 13'sd 4033) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14597) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11871) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27678) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25307) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13455) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29640) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11425) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16571) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9368) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20384) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1831) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18677) * $signed(input_fmap_107[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3088) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11607) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_112[7:0]) +
	( 10'sd 394) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6062) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21661) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30558) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11992) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3371) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25107) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26740) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 15'sd 14883) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29493) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1698) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31028) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5698) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25555) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26192) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26870) * $signed(input_fmap_9[7:0]) +
	( 11'sd 745) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5871) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25286) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27365) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21993) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12233) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9005) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17704) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1849) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23640) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18334) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6861) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17970) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19318) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5293) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21210) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23918) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16933) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2456) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17547) * $signed(input_fmap_39[7:0]) +
	( 9'sd 154) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31723) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16455) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1122) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7742) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29626) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4184) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6113) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5151) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21972) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27970) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15428) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27776) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19802) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26612) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23634) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15213) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31201) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6162) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10797) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18639) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16299) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32534) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_72[7:0]) +
	( 13'sd 4018) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14638) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_75[7:0]) +
	( 10'sd 264) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12401) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25348) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1412) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6705) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21240) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_83[7:0]) +
	( 10'sd 291) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31190) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3398) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9788) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7735) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21701) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31640) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9400) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7669) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4216) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15348) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14305) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15202) * $signed(input_fmap_101[7:0]) +
	( 9'sd 139) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2749) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16363) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24344) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1603) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14874) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7694) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6415) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25576) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18294) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10569) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17059) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1868) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15185) * $signed(input_fmap_123[7:0]) +
	( 8'sd 87) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28621) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15680) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 14'sd 4302) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30462) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29562) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17128) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16476) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16629) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28246) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28388) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32317) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21630) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3314) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22039) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11293) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16127) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28466) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5823) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1751) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25453) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12839) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10947) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18282) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31456) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15794) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11314) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24514) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23425) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30187) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19669) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21885) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2277) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29055) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10774) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23048) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6358) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28137) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5276) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1969) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13608) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23535) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9112) * $signed(input_fmap_62[7:0]) +
	( 10'sd 313) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6997) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3360) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24853) * $signed(input_fmap_66[7:0]) +
	( 9'sd 240) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29397) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31988) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14140) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6729) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29477) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10451) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19201) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10128) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4747) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14683) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29747) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6949) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13348) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21161) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3563) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26558) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7036) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14441) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26700) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18973) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15087) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23587) * $signed(input_fmap_101[7:0]) +
	( 10'sd 316) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32274) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16597) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16334) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4897) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23159) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10589) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30649) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24034) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3895) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18796) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29848) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8037) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29852) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28186) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12510) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 16'sd 20727) * $signed(input_fmap_0[7:0]) +
	( 11'sd 829) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12648) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31458) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6098) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4964) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17319) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17096) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11554) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25856) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1378) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16031) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12864) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27007) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20401) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24224) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1671) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12517) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7791) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2342) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16369) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24760) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24444) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25945) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22582) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16549) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13406) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24904) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3627) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18031) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11670) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18171) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15384) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_56[7:0]) +
	( 10'sd 494) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10363) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31599) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16092) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7843) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30568) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5929) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8672) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12601) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13255) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9711) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17157) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9114) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25847) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30036) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11025) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18021) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9180) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31072) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30718) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28485) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_85[7:0]) +
	( 11'sd 925) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23687) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16190) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15254) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26361) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28195) * $signed(input_fmap_91[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_93[7:0]) +
	( 11'sd 709) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3774) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29577) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27590) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22710) * $signed(input_fmap_106[7:0]) +
	( 10'sd 377) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24607) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27195) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11081) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16382) * $signed(input_fmap_114[7:0]) +
	( 13'sd 4052) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15379) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11999) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5823) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13734) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31050) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 16'sd 19332) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17336) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3887) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25079) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27421) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11927) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11856) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8016) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20953) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22013) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15463) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25151) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7423) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11077) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31909) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13078) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15204) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19609) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32530) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2411) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29256) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28002) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_35[7:0]) +
	( 11'sd 586) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10528) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21953) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22460) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27712) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18710) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5793) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16810) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27023) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13511) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23777) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10215) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7903) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14062) * $signed(input_fmap_58[7:0]) +
	( 10'sd 375) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20499) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17050) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5134) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12617) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20092) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32347) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24810) * $signed(input_fmap_70[7:0]) +
	( 10'sd 453) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26941) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6082) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21831) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6276) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19407) * $signed(input_fmap_78[7:0]) +
	( 11'sd 693) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22560) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5716) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31780) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9187) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7288) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17758) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14087) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_90[7:0]) +
	( 11'sd 981) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_92[7:0]) +
	( 10'sd 365) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20236) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10588) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19765) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25027) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15545) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3550) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16320) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10506) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13095) * $signed(input_fmap_103[7:0]) +
	( 7'sd 62) * $signed(input_fmap_104[7:0]) +
	( 11'sd 977) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6550) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17930) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23294) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15490) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9840) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2843) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10002) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24983) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22282) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30584) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1636) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9495) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32011) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 16'sd 30504) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18237) * $signed(input_fmap_2[7:0]) +
	( 10'sd 402) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18190) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19954) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28104) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28938) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10521) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26287) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17294) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15528) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7486) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29471) * $signed(input_fmap_15[7:0]) +
	( 11'sd 999) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9351) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20190) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4253) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2050) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23674) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16960) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7770) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29817) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16953) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4954) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4378) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5647) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29232) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13270) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8862) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30427) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15009) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19143) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32079) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23301) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18659) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14907) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30561) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16919) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9350) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21266) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10052) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5163) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27572) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10585) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26615) * $signed(input_fmap_70[7:0]) +
	( 11'sd 614) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27178) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25654) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3651) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1585) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12016) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22608) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32001) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7864) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28784) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24794) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15683) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17522) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8242) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2832) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32483) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12282) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8350) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17179) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31470) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5504) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3415) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3056) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7368) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19115) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22026) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3094) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29331) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23912) * $signed(input_fmap_113[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13796) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6674) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30177) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12067) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4182) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21742) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27960) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10516) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 16'sd 19639) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15941) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30919) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31525) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13044) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28930) * $signed(input_fmap_11[7:0]) +
	( 11'sd 677) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28670) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27244) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18057) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8913) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20203) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14059) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31249) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31469) * $signed(input_fmap_24[7:0]) +
	( 10'sd 487) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10879) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32553) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3913) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25707) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18167) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18627) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10010) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13658) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18469) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11624) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22582) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15693) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3408) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15521) * $signed(input_fmap_44[7:0]) +
	( 7'sd 50) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11231) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1801) * $signed(input_fmap_47[7:0]) +
	( 11'sd 816) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12553) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20704) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1261) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13189) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27989) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7922) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23440) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10329) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15985) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12340) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19744) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24794) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26893) * $signed(input_fmap_67[7:0]) +
	( 11'sd 902) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2673) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16199) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20322) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22655) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5130) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23783) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20004) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31271) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14662) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20383) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25938) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27366) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15598) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20270) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9941) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5934) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22330) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1209) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6626) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27417) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18453) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4900) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9384) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24097) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3841) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24970) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19521) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28028) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29411) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20356) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24225) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12919) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3300) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3250) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15081) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10521) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2849) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 16'sd 21751) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4326) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14409) * $signed(input_fmap_2[7:0]) +
	( 11'sd 551) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10597) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19492) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14670) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22398) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8451) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10953) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18502) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2648) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30058) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27513) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23896) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25597) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25006) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20419) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31680) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1946) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6407) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5298) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5483) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24784) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24801) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31212) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7326) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32022) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10885) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10984) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12461) * $signed(input_fmap_45[7:0]) +
	( 11'sd 614) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13934) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12670) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25507) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1265) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16672) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24165) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24940) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20648) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12578) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9291) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27767) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1151) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1992) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28496) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3216) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10776) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12641) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25088) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26260) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27216) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31776) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2130) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12959) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22844) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11132) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27424) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32152) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7105) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8831) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4204) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16376) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18878) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9628) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25982) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15960) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24215) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_101[7:0]) +
	( 11'sd 513) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31067) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27604) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12388) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10589) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6453) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8712) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19559) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10238) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4547) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19233) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10806) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_117[7:0]) +
	( 8'sd 109) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11859) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9936) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14711) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 15'sd 14451) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5217) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14613) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5255) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2170) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22562) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5776) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31986) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9771) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30381) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31004) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32549) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24245) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22034) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2454) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22269) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3810) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32260) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16299) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7765) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1593) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13415) * $signed(input_fmap_33[7:0]) +
	( 11'sd 541) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11309) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6032) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21654) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3690) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30807) * $signed(input_fmap_43[7:0]) +
	( 9'sd 141) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29703) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18948) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19961) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26087) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18207) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22520) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25700) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17604) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8045) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31215) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3175) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2306) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9802) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25549) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29465) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1995) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20116) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31355) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12394) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4456) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32011) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27381) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3785) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5104) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21251) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25137) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2894) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30769) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7330) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11899) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23594) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6658) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21627) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7734) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20834) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3280) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23466) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5443) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20039) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3630) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12510) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5083) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22753) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22775) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22841) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18586) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16248) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11349) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24346) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17845) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17729) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31319) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6072) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 14'sd 7052) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10240) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16224) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32262) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12253) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11189) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9026) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32416) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29663) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16576) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11798) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_20[7:0]) +
	( 13'sd 4014) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4689) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28539) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2762) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7924) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23711) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16952) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14144) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27894) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28172) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13467) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27019) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23953) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21028) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10446) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2538) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31650) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22949) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26745) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2065) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23287) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13627) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25909) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20567) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20943) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12556) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27360) * $signed(input_fmap_61[7:0]) +
	( 12'sd 2027) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9241) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20519) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29024) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24923) * $signed(input_fmap_72[7:0]) +
	( 10'sd 281) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4248) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8774) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28993) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1389) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32653) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24695) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1791) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22380) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27241) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8780) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15772) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29396) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28283) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5943) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1295) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31426) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28346) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29968) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8509) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18325) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13765) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7827) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18982) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15828) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9712) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22217) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19331) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25458) * $signed(input_fmap_113[7:0]) +
	( 11'sd 819) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14425) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 16'sd 17419) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1380) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29609) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6148) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21671) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8606) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4143) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27887) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32285) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24296) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23889) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24185) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25574) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19526) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25374) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23357) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4517) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22445) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5009) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1179) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7422) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31521) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27698) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17000) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2944) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28233) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27600) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17149) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28205) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17192) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28712) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3338) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31886) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20069) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21207) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20008) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28378) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1312) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22054) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31768) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18493) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2088) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13477) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3277) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27165) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8561) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24467) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23597) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25227) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25459) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14551) * $signed(input_fmap_76[7:0]) +
	( 9'sd 134) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28901) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11894) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26671) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12189) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30917) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25809) * $signed(input_fmap_86[7:0]) +
	( 3'sd 3) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30665) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30655) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11021) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22081) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14387) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11434) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31097) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25599) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25190) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15367) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17042) * $signed(input_fmap_106[7:0]) +
	( 8'sd 112) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27284) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8909) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8535) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28755) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_116[7:0]) +
	( 12'sd 2037) * $signed(input_fmap_117[7:0]) +
	( 10'sd 373) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19467) * $signed(input_fmap_119[7:0]) +
	( 11'sd 1022) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21992) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14259) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18116) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17907) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3647) * $signed(input_fmap_125[7:0]) +
	( 11'sd 970) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_127[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 12'd1537;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 16'd18702;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 16'd20624;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 15'd9373;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 13'd3158;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 15'd8804;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 16'd26181;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 15'd11456;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 15'd9150;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 16'd29033;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 16'd20346;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 14'd6119;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 16'd31466;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 16'd23933;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 13'd2124;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 16'd27688;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 8'd64;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 16'd24268;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 16'd25926;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 14'd5535;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 16'd16959;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 16'd27651;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 15'd11401;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 14'd7101;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 16'd32585;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 12'd1231;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 15'd12902;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 14'd5033;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 14'd5483;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 14'd5373;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 16'd19606;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 15'd12854;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 11'd734;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 15'd12838;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 16'd31238;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 14'd6588;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 12'd1556;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 16'd21692;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 16'd22679;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 16'd17386;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 16'd18837;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 13'd2466;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 16'd23457;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 16'd28617;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 14'd5585;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 15'd10025;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 14'd6897;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 16'd30482;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 15'd16167;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 16'd19125;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 15'd12637;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 15'd15055;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 15'd16288;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 13'd2407;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 16'd17503;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 15'd10252;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 10'd436;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 16'd26109;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 8'd104;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 16'd28086;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 15'd12953;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 15'd8634;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 16'd22347;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 16'd25920;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 14'd4947;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 15'd9854;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 16'd26673;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 14'd4860;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 16'd31592;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 13'd2503;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 15'd12440;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 15'd16019;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 15'd11243;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 16'd17332;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 14'd4400;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 16'd31780;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 15'd12373;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 10'd433;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 16'd25263;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 16'd17473;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 16'd29203;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 12'd1861;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 16'd18294;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 16'd27817;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 16'd20327;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 16'd22219;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 15'd14084;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 15'd9231;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 15'd14213;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 16'd19744;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 16'd25415;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 16'd27280;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 15'd10924;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 16'd28773;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 16'd29402;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 15'd13734;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 16'd17346;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 16'd32043;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 16'd22308;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 15'd9256;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 14'd4836;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 14'd7864;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 16'd32075;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 16'd30940;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 16'd27922;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 15'd10923;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 14'd6739;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 16'd27118;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 16'd22596;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 14'd4227;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 16'd25824;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 12'd1771;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 15'd10195;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 16'd28294;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 16'd25103;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 15'd15530;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 15'd10781;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 15'd11099;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 16'd22909;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 16'd17656;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 15'd8904;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 12'd1528;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 16'd31515;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 12'd1816;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 15'd15203;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 14'd5103;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 15'd13406;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 14'd6612;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[21:15]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[21:15]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[21:15]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[21:15]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[21:15]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[21:15]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[21:15]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[21:15]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[21:15]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[21:15]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[21:15]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[21:15]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[21:15]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[21:15]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[21:15]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[21:15]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[21:15]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[21:15]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[21:15]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[21:15]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[21:15]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[21:15]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[21:15]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[21:15]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[21:15]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[21:15]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[21:15]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[21:15]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[21:15]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[21:15]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[21:15]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[21:15]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[21:15]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[21:15]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[21:15]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[21:15]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[21:15]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[21:15]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[21:15]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[21:15]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[21:15]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[21:15]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[21:15]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[21:15]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[21:15]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[21:15]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[21:15]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[21:15]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[21:15]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[21:15]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[21:15]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[21:15]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[21:15]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[21:15]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[21:15]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[21:15]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[21:15]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[21:15]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[21:15]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[21:15]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[21:15]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[21:15]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[21:15]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[21:15]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[21:15]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[21:15]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[21:15]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[21:15]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[21:15]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[21:15]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[21:15]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[21:15]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[21:15]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[21:15]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[21:15]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[21:15]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[21:15]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[21:15]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[21:15]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[21:15]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[21:15]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[21:15]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[21:15]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[21:15]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[21:15]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[21:15]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[21:15]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[21:15]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[21:15]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[21:15]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[21:15]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[21:15]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[21:15]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[21:15]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[21:15]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[21:15]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[21:15]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[21:15]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[21:15]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[21:15]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[21:15]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[21:15]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[21:15]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[21:15]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[21:15]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[21:15]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[21:15]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[21:15]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[21:15]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[21:15]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[21:15]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[21:15]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[21:15]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[21:15]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[21:15]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[21:15]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[21:15]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[21:15]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[21:15]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[21:15]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[21:15]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[21:15]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[21:15]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[21:15]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[21:15]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[21:15]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[21:15]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[21:15]}} :'d6) : '0;

assign output_act = {
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
