module conv10_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [1024-1:0] input_act,
    output logic [1024-1:0] output_act,
    output logic ready
);

logic [1024-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 16'sd 27910) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16257) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12833) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16378) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21828) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26975) * $signed(input_fmap_5[7:0]) +
	( 11'sd 532) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23334) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23418) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_10[7:0]) +
	( 9'sd 190) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32504) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24620) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13343) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5561) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17758) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1626) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3090) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21273) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3450) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9147) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26292) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8355) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31423) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9866) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28306) * $signed(input_fmap_34[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21583) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22166) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29605) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20031) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22203) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3763) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27376) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26764) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8344) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11882) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16559) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12169) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1937) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21911) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6738) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18518) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6715) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4609) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29652) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5367) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24785) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7478) * $signed(input_fmap_66[7:0]) +
	( 13'sd 4091) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20384) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13349) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20578) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27228) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14194) * $signed(input_fmap_75[7:0]) +
	( 5'sd 11) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18997) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23713) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5067) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19035) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18722) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18764) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3565) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19922) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9243) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_90[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15212) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_93[7:0]) +
	( 11'sd 864) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13021) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21599) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27593) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2454) * $signed(input_fmap_100[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17691) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9487) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30037) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8527) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12569) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15017) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28597) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16278) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8299) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15448) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16966) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22247) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2858) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15177) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29858) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27827) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 16'sd 22959) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27558) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7938) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18621) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4324) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30415) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21153) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24740) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18288) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15383) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9731) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24940) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13872) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14262) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1526) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22244) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32039) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27589) * $signed(input_fmap_31[7:0]) +
	( 11'sd 859) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19934) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16134) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32211) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18560) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21857) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22287) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12490) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27919) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25298) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32716) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25390) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13680) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17928) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27928) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12301) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6972) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2269) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26787) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11989) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8754) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28904) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16664) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22725) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31482) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_68[7:0]) +
	( 11'sd 904) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2478) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21492) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9952) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26725) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5795) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30361) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8437) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18574) * $signed(input_fmap_85[7:0]) +
	( 11'sd 708) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29986) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24665) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16326) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31618) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2471) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7088) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19997) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16312) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21158) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21477) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18425) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30823) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2192) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14910) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22116) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17930) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16123) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27008) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10236) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6407) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28259) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11085) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19390) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11950) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1563) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11394) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22088) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3863) * $signed(input_fmap_126[7:0]) +
	( 11'sd 685) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 16'sd 22772) * $signed(input_fmap_0[7:0]) +
	( 14'sd 8187) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20489) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6229) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9297) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19872) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5186) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26524) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31299) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9537) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31150) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18266) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25215) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5760) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5935) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26489) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_22[7:0]) +
	( 11'sd 800) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7734) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5562) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4184) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15329) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19249) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14119) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27403) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3710) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32183) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8563) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11060) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26168) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16508) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31147) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24077) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21775) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32615) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18049) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2760) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23002) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15710) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32256) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28463) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24396) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21281) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5149) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19298) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1869) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30099) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16651) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23599) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16155) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10555) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_87[7:0]) +
	( 11'sd 732) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12997) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30383) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7067) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17810) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22480) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14146) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9211) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23199) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11517) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9273) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31521) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14209) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23344) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13919) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27798) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17955) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11957) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20692) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31001) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30694) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30692) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9384) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5356) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4844) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11728) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21560) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2695) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21238) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 16'sd 22846) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21657) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16955) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_4[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5743) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_7[7:0]) +
	( 11'sd 604) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7786) * $signed(input_fmap_9[7:0]) +
	( 11'sd 896) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4542) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15384) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16131) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19220) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12462) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3690) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12634) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20166) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25621) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10947) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14162) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20404) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9063) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31167) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29766) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20798) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6086) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30509) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4432) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26205) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4825) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13305) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19322) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5299) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_44[7:0]) +
	( 13'sd 4006) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28060) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31852) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22127) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31705) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11698) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5531) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16795) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27403) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1476) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13490) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3531) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32740) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25474) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3380) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7951) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9556) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8500) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21463) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2157) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25119) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15397) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4466) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31537) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8924) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10860) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30663) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8866) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24130) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9712) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23343) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16019) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28033) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27712) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9795) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17433) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5460) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1030) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_109[7:0]) +
	( 11'sd 750) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10422) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17262) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21206) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13265) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22046) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14508) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1798) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6430) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 15'sd 11864) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10503) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4588) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18445) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14360) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_6[7:0]) +
	( 13'sd 4041) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27687) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15097) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31139) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12496) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1780) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7683) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13838) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11348) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7095) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26973) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2077) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3184) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12351) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30356) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7799) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23778) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13332) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11176) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28892) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17302) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12114) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28471) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5617) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3174) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15970) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8637) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21624) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16010) * $signed(input_fmap_50[7:0]) +
	( 10'sd 472) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29498) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23587) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17867) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11200) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6532) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19180) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20059) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8525) * $signed(input_fmap_70[7:0]) +
	( 13'sd 4068) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7616) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20725) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25634) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22000) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9484) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31870) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18820) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_89[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31630) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26233) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14118) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17126) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18068) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23247) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9332) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11111) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6444) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25746) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5366) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16622) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16516) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25138) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16482) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6414) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30575) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30837) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9341) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28883) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27757) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 13'sd 2086) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7906) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19509) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23785) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11995) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24018) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_8[7:0]) +
	( 8'sd 100) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16424) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_12[7:0]) +
	( 11'sd 658) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23125) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2557) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21960) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21060) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4926) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28412) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6388) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9517) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2354) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29553) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3809) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1365) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2669) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23373) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30266) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18394) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19330) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8933) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1206) * $signed(input_fmap_45[7:0]) +
	( 13'sd 4005) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1444) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27607) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27509) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25427) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22782) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26769) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9173) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14989) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29277) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5030) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3937) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19236) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15106) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1426) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26102) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1675) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23666) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8011) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6739) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9610) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31194) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23211) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25610) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12775) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25222) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14114) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31450) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2688) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6915) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5474) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27291) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26184) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22480) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28572) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25936) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31259) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16988) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14908) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5882) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12789) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26340) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30905) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4432) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5364) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21676) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13170) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21560) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10519) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15728) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29229) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18188) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16631) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 16'sd 25501) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30278) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3208) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26596) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4345) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14524) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7876) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21775) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23446) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24083) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21896) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18655) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29525) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21356) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19024) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8275) * $signed(input_fmap_20[7:0]) +
	( 14'sd 8021) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2942) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6040) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11939) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9960) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5741) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26029) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15321) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30911) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24193) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19021) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7013) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17442) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2793) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20098) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16555) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24130) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30260) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32692) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26297) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14249) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28721) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12883) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5033) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13790) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16119) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27811) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25009) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29841) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5665) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22850) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25831) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13132) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13786) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7325) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24754) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15062) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2335) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13982) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15956) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18995) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11839) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12759) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14808) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18754) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5483) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6246) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24427) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8291) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31790) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9144) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30087) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16167) * $signed(input_fmap_84[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26889) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18476) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1039) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26803) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19662) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13598) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29609) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6252) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26150) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19534) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27543) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30386) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22754) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19160) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4600) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7735) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31068) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7910) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11937) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30618) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13052) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20846) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25609) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22189) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15454) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 16'sd 29041) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12747) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4282) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8278) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14642) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2071) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22658) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1649) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1458) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26909) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5230) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25511) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20625) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6931) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5378) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3440) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13507) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27807) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32609) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29257) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3676) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2218) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7583) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26024) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15172) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31441) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21126) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30609) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15763) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23155) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23960) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20228) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4290) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1805) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11673) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10879) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28055) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6318) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5921) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10546) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27782) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27187) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27794) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11674) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10345) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8086) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13926) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29587) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21937) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1262) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7048) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16152) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21017) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4739) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6936) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16050) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30511) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27157) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8958) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14448) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31841) * $signed(input_fmap_96[7:0]) +
	( 12'sd 2012) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15816) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17124) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8977) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26290) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20072) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3391) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14317) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32122) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9189) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9772) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27026) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18534) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11697) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16834) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14670) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20702) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30605) * $signed(input_fmap_123[7:0]) +
	( 11'sd 998) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14078) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 14'sd 7397) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22806) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30813) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1976) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32590) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11899) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30538) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11711) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17939) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10685) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19963) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16250) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19491) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26116) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20784) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7198) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27548) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27385) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21967) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6866) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24819) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25556) * $signed(input_fmap_36[7:0]) +
	( 11'sd 604) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29612) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13653) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3419) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4749) * $signed(input_fmap_42[7:0]) +
	( 8'sd 91) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31499) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23583) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25240) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9524) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12408) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29619) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30085) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1505) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16466) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5517) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23764) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1530) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9068) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2352) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25477) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22466) * $signed(input_fmap_67[7:0]) +
	( 8'sd 98) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24980) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5767) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5809) * $signed(input_fmap_73[7:0]) +
	( 10'sd 366) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1985) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21978) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28310) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11081) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24529) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31953) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19704) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22731) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15911) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31052) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1797) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14790) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17523) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5120) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27391) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27360) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16788) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6640) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25290) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27619) * $signed(input_fmap_102[7:0]) +
	( 11'sd 540) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19745) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11678) * $signed(input_fmap_106[7:0]) +
	( 8'sd 70) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16752) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1765) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15679) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21727) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3074) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12087) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18726) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7341) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21161) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27507) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6075) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 16'sd 25885) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7879) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5716) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20711) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29244) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5714) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7643) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28117) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17872) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22037) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25831) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10050) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14036) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26180) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17445) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7021) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14209) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24725) * $signed(input_fmap_19[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26229) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30308) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8410) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4369) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17204) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14913) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29217) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13511) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4434) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2681) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25174) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31844) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23738) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25830) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9595) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26795) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3755) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5664) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19076) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14287) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11088) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30152) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27698) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29228) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19856) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9772) * $signed(input_fmap_54[7:0]) +
	( 11'sd 756) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12546) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15700) * $signed(input_fmap_57[7:0]) +
	( 9'sd 158) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3934) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8151) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32692) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26920) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25347) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22790) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7826) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13519) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3601) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17195) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12977) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30621) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6564) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10789) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10305) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25234) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22897) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2515) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27162) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14467) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4124) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16495) * $signed(input_fmap_88[7:0]) +
	( 8'sd 84) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3708) * $signed(input_fmap_92[7:0]) +
	( 11'sd 1000) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32515) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23061) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20198) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13958) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4978) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5285) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14375) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13311) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30349) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26418) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16917) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22065) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15972) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15556) * $signed(input_fmap_117[7:0]) +
	( 9'sd 253) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14588) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23023) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20343) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6534) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11368) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30581) * $signed(input_fmap_125[7:0]) +
	( 9'sd 236) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27335) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 16'sd 16880) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14997) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13694) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22912) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27950) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2167) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1431) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22161) * $signed(input_fmap_10[7:0]) +
	( 12'sd 2023) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29700) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12299) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24407) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8320) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1029) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32308) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23025) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11160) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6804) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31987) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32665) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17402) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14926) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10182) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10395) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22453) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24962) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28913) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2676) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30939) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1901) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15199) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21536) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4880) * $signed(input_fmap_47[7:0]) +
	( 11'sd 935) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23427) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_52[7:0]) +
	( 11'sd 900) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19198) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18442) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23796) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30588) * $signed(input_fmap_64[7:0]) +
	( 11'sd 644) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7649) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16083) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17426) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15652) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15926) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16298) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29826) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21158) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1475) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12853) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2353) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25997) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13760) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4815) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_84[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1955) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32678) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21757) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1748) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8213) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20713) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13998) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4953) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2971) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21201) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31505) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3985) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22391) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10839) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25679) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23756) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21222) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26258) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29944) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3990) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20202) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27029) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 15'sd 15954) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18200) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25057) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15655) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19977) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2704) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30884) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13635) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15912) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22363) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16376) * $signed(input_fmap_16[7:0]) +
	( 11'sd 828) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17760) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20211) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20971) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11147) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32305) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6649) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14439) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_29[7:0]) +
	( 11'sd 828) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11781) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22850) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17757) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6606) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10991) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26409) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19224) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9858) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12634) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28443) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14227) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22832) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11285) * $signed(input_fmap_49[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2816) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27133) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17498) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29287) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32680) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23107) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13365) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25372) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28698) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32686) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23162) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6770) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9572) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18396) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22283) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3407) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19891) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31467) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17328) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27809) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14678) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3146) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3966) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7926) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21718) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25676) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15375) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32394) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21484) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17677) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24230) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10240) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9960) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21069) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6596) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27580) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1370) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7001) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25020) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31157) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17757) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26311) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19784) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 15'sd 10101) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7709) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18300) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25443) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8880) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9920) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17809) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27125) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17212) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14707) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8362) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32194) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17902) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2946) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9448) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11271) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10522) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13354) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20801) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5725) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31568) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14331) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23771) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6190) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12009) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30435) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7976) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27270) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2959) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8381) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30995) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2241) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1573) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23361) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13700) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9275) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18643) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24280) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3492) * $signed(input_fmap_58[7:0]) +
	( 10'sd 492) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4505) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17874) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2322) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26556) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13372) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12025) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11937) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14594) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9560) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16478) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2781) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12805) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28241) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16339) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9147) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32636) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15276) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28446) * $signed(input_fmap_90[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30736) * $signed(input_fmap_93[7:0]) +
	( 14'sd 8129) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17069) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3849) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26592) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18798) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19577) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27966) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28017) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4125) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30561) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9658) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4630) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25763) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9194) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18704) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21900) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15384) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23458) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11293) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20999) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27679) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 16'sd 19927) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10347) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28156) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25336) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4738) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13978) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29497) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12684) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15685) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19665) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5192) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3370) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16966) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2318) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28896) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31078) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22691) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22119) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10654) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9644) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29990) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30271) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28711) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16666) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23433) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_40[7:0]) +
	( 11'sd 1007) * $signed(input_fmap_41[7:0]) +
	( 11'sd 684) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24916) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22518) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8486) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13928) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12462) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2625) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29513) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30411) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13114) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7636) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11108) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28629) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24054) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29291) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23023) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3574) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6400) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32683) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2654) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7663) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32759) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8943) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17018) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29317) * $signed(input_fmap_80[7:0]) +
	( 13'sd 4086) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19007) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9247) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16830) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12214) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30012) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13581) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5067) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22496) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11915) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21342) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13022) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31471) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31138) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7703) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10302) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28026) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8113) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27402) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30921) * $signed(input_fmap_113[7:0]) +
	( 8'sd 110) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14124) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23822) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5606) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11318) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20807) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1638) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17925) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_125[7:0]) +
	( 9'sd 134) * $signed(input_fmap_126[7:0]) +
	( 7'sd 62) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 16'sd 18852) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23677) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8953) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10101) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32107) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28896) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23988) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25938) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19334) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23298) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3058) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13804) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22318) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13337) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6918) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1836) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1290) * $signed(input_fmap_24[7:0]) +
	( 5'sd 8) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26144) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31157) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31872) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14808) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18898) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22760) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27455) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30056) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19942) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16152) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20802) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10819) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7682) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18410) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3848) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3229) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10163) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11951) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7365) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28740) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22599) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19408) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16917) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11742) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18261) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25594) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31237) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14808) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27571) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12149) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15848) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13383) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4370) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20182) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16666) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24111) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26414) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15831) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9043) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20863) * $signed(input_fmap_91[7:0]) +
	( 10'sd 413) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13804) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28348) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15619) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17594) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11136) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11288) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27298) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29377) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29198) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2946) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14252) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2854) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8443) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32044) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32455) * $signed(input_fmap_117[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18929) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4416) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6390) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21982) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17809) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 13'sd 2668) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32675) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29480) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28432) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19797) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11539) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31281) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22411) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26584) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_12[7:0]) +
	( 8'sd 124) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6709) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15289) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15508) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19431) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31974) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2878) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10319) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19291) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19160) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10128) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27464) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5345) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26684) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11647) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30395) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20259) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27981) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27044) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23993) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5667) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11434) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11214) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6964) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32717) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29327) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25019) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23049) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15343) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2891) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14224) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22968) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28018) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28949) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2948) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4323) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1633) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11554) * $signed(input_fmap_76[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7351) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25930) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15061) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25094) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29797) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9943) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19781) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32229) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12783) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10104) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4587) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18208) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25746) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4409) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1186) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2797) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3850) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31922) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3830) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6000) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8883) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23791) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16648) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7703) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1461) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19258) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3167) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2481) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19557) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20900) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6752) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20409) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19751) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7414) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26302) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 14'sd 7348) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6515) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10947) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29249) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10464) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9701) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11535) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22456) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30156) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10713) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15044) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24638) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2325) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19883) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23519) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1730) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11025) * $signed(input_fmap_22[7:0]) +
	( 10'sd 462) * $signed(input_fmap_23[7:0]) +
	( 10'sd 482) * $signed(input_fmap_24[7:0]) +
	( 10'sd 364) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_26[7:0]) +
	( 8'sd 103) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25379) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26414) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21679) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19695) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14469) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30377) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7209) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5058) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19690) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2783) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17724) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9910) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20554) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4354) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2128) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5786) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17071) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14303) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2408) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14769) * $signed(input_fmap_61[7:0]) +
	( 14'sd 8076) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_63[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5041) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23725) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18973) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18414) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8395) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28588) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_76[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28901) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6141) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23211) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13306) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31273) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12098) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28025) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4826) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12481) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6504) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5597) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7246) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23763) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9805) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29402) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30454) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18735) * $signed(input_fmap_102[7:0]) +
	( 10'sd 422) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28052) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3907) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25876) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31700) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14986) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27039) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31558) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30845) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4560) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7733) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24556) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28524) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31388) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30998) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25840) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21744) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10721) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 14'sd 5412) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11352) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11674) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23821) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1811) * $signed(input_fmap_5[7:0]) +
	( 12'sd 2027) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12746) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14737) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3514) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23382) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27812) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23366) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7800) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1960) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15262) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4457) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16447) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28570) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30432) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12386) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7142) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23255) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9696) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6652) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28016) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17265) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7502) * $signed(input_fmap_43[7:0]) +
	( 9'sd 217) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9964) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18432) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8888) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23390) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27848) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12697) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28842) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22511) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16410) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19000) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29180) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8401) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24772) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9896) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11356) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9536) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24699) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21098) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17090) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12915) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10891) * $signed(input_fmap_78[7:0]) +
	( 11'sd 977) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19976) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31371) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23665) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14908) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11942) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22915) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5810) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10991) * $signed(input_fmap_89[7:0]) +
	( 10'sd 267) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19700) * $signed(input_fmap_91[7:0]) +
	( 11'sd 741) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12138) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31321) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_95[7:0]) +
	( 11'sd 689) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_99[7:0]) +
	( 12'sd 2011) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4315) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17294) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28566) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22664) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17603) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13696) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10519) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28065) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25015) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2446) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_120[7:0]) +
	( 10'sd 459) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16533) * $signed(input_fmap_122[7:0]) +
	( 10'sd 395) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16325) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19380) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 16'sd 30259) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27165) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20576) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7002) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8512) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26079) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28325) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20956) * $signed(input_fmap_12[7:0]) +
	( 11'sd 786) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5029) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20305) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2860) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16606) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10581) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25354) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16454) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6038) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14543) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11029) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17984) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3594) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16196) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31366) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24865) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23593) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29835) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28406) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15781) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31691) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3738) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9942) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8902) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7315) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20638) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19502) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5567) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18241) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27494) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2671) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3322) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30166) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1796) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_65[7:0]) +
	( 10'sd 351) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30572) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6141) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12496) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13406) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20100) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1678) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28849) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11441) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32258) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2055) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9232) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30029) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6723) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28202) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18472) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15019) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4229) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12096) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6957) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22251) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26876) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22175) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18362) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11856) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32354) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2263) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29903) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18585) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16797) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1871) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22334) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3122) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18695) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_123[7:0]) +
	( 10'sd 277) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12867) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4182) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 15'sd 11027) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12143) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12299) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17440) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18628) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13565) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12821) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16344) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9562) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25931) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10406) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5736) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26740) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3858) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7005) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12634) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22711) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16922) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29421) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29618) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28542) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18230) * $signed(input_fmap_33[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21539) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3534) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26744) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6199) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17517) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27732) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7855) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24359) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23656) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27753) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13366) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29311) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2162) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9578) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30537) * $signed(input_fmap_55[7:0]) +
	( 11'sd 722) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8309) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14067) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12387) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_61[7:0]) +
	( 13'sd 4049) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14027) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12825) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11556) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19706) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18190) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7916) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10809) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2377) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32359) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28925) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13633) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30731) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24905) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14634) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13886) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20731) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31165) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25774) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28295) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14202) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7874) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23137) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5148) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7296) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21348) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2279) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17659) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9660) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23577) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12345) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28857) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20655) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5411) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32578) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15115) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20388) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12080) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5125) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15181) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6621) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 16'sd 20552) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21324) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19166) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5865) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2715) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3371) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24970) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29199) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30709) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7380) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11295) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28249) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20508) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1966) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16657) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23466) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10999) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32357) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12346) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32027) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25781) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15488) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13936) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14736) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20576) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31341) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24830) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19479) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1610) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10136) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22038) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20659) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22659) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22960) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2348) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22388) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_58[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5199) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8723) * $signed(input_fmap_62[7:0]) +
	( 11'sd 854) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22956) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6121) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28583) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15383) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15831) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27963) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6101) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15787) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25459) * $signed(input_fmap_75[7:0]) +
	( 11'sd 572) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22696) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22898) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8285) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9288) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19787) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27335) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12891) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26342) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2672) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30617) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16406) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24243) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7948) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32346) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5096) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11822) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17851) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8282) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15508) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32739) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26916) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2264) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5282) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7026) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19629) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31528) * $signed(input_fmap_114[7:0]) +
	( 10'sd 492) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24065) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25159) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12305) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20945) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24806) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24584) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13916) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6023) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30195) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 15'sd 9167) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29497) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6498) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16935) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6290) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28469) * $signed(input_fmap_8[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23265) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30886) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6898) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23533) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19267) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13522) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21801) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5536) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7324) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8734) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7923) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19418) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1428) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_33[7:0]) +
	( 10'sd 400) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28986) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16192) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4451) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19531) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26031) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29673) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14683) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14641) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7737) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6461) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17813) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16646) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21052) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17959) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23199) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11453) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19329) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4755) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12487) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27801) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_65[7:0]) +
	( 11'sd 850) * $signed(input_fmap_66[7:0]) +
	( 10'sd 471) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24978) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_70[7:0]) +
	( 9'sd 220) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19151) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21545) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27963) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9134) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1437) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11480) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19884) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20957) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14752) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14202) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_86[7:0]) +
	( 11'sd 611) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5819) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7009) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21967) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2765) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16477) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11510) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8909) * $signed(input_fmap_98[7:0]) +
	( 8'sd 120) * $signed(input_fmap_99[7:0]) +
	( 13'sd 4010) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13195) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2365) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31362) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1463) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29887) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22545) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1584) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24510) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7951) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29459) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15324) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2959) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2411) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10209) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32755) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 15'sd 11035) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15980) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7106) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4597) * $signed(input_fmap_4[7:0]) +
	( 11'sd 928) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9568) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10020) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2646) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28394) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26056) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25405) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22289) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10536) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9311) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20682) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22530) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16556) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19164) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10209) * $signed(input_fmap_25[7:0]) +
	( 10'sd 508) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7920) * $signed(input_fmap_27[7:0]) +
	( 11'sd 634) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24441) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11286) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12182) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14258) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18874) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2384) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14352) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11155) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17553) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25862) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11661) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23645) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10481) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3523) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4822) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16861) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5980) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31530) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12842) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13319) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22268) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13846) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27578) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5369) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14569) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11940) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18933) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6723) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28029) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7718) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26631) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18631) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7195) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29165) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29340) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17436) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_84[7:0]) +
	( 9'sd 239) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3921) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12428) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11018) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4763) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11081) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10731) * $signed(input_fmap_95[7:0]) +
	( 10'sd 361) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23554) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25058) * $signed(input_fmap_101[7:0]) +
	( 11'sd 906) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20735) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17750) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16534) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29711) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32032) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_110[7:0]) +
	( 11'sd 864) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15780) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25080) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1826) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27474) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12341) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12404) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8067) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11706) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_125[7:0]) +
	( 9'sd 182) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18763) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 15'sd 9567) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19695) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10706) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31460) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26460) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15505) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32635) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14409) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_11[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2092) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1044) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7144) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18918) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31076) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22565) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17357) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20846) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11091) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13132) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1142) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32251) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7528) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16304) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30281) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18354) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14178) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12085) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5441) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19035) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29551) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25220) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5159) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26687) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4305) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24415) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3057) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23172) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28675) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23462) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5553) * $signed(input_fmap_55[7:0]) +
	( 15'sd 16180) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9063) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16344) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2207) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3088) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14704) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27121) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7027) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28921) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12314) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1024) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22926) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2679) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15075) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22821) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27195) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16282) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18209) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11269) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1230) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12553) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19316) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18767) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5726) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12143) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29625) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11872) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11057) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6409) * $signed(input_fmap_99[7:0]) +
	( 14'sd 8154) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16070) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21061) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17487) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22317) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27563) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14024) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18052) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3476) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25029) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6134) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23832) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22578) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16830) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10670) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12078) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32332) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31253) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 14'sd 5130) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26277) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27141) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28453) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8831) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30567) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25175) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32299) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20218) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_18[7:0]) +
	( 9'sd 205) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3752) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15394) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17582) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10673) * $signed(input_fmap_25[7:0]) +
	( 13'sd 4042) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6567) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25569) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9816) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28870) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10842) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12759) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15193) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22883) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6614) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20031) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21315) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15651) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24605) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16587) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30089) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22935) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24348) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22978) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19589) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27110) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25404) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8249) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19190) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_77[7:0]) +
	( 11'sd 624) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24950) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26853) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4857) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2785) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1336) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10677) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12172) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29328) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18493) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8955) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7252) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15775) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6219) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14965) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32366) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23301) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2308) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9576) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23077) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14208) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17420) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32594) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18959) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3335) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9182) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5072) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11703) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11754) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20950) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11933) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10754) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19828) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28552) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18056) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27061) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2837) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3561) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26883) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26091) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 16'sd 17290) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3554) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12520) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21883) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4670) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24423) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25538) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9760) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26700) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18352) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10269) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6381) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29017) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26211) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11603) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19382) * $signed(input_fmap_30[7:0]) +
	( 10'sd 388) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5075) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2166) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22701) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6725) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20994) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16580) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18142) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18971) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15355) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20793) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15621) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27820) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31869) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30634) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17596) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12439) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29554) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25177) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1604) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31058) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5835) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13936) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12112) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22338) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32400) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27663) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12462) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18959) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3532) * $signed(input_fmap_80[7:0]) +
	( 8'sd 110) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22795) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26874) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5504) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27496) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11454) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11755) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4208) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3060) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30510) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2353) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_95[7:0]) +
	( 13'sd 4031) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14296) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26622) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16472) * $signed(input_fmap_99[7:0]) +
	( 9'sd 197) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_101[7:0]) +
	( 9'sd 187) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25630) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8597) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27355) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5353) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18099) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26811) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29770) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21935) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8469) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2270) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19861) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_121[7:0]) +
	( 8'sd 106) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1661) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21733) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_125[7:0]) +
	( 9'sd 222) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26197) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 14'sd 6306) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29378) * $signed(input_fmap_1[7:0]) +
	( 10'sd 492) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14336) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16334) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25073) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1142) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9025) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12333) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23647) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21919) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31421) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12153) * $signed(input_fmap_24[7:0]) +
	( 10'sd 486) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12913) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14620) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27533) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31061) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11335) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25624) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22731) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8915) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19813) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27969) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31397) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19797) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28751) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6923) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19599) * $signed(input_fmap_49[7:0]) +
	( 10'sd 284) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5834) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14967) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27565) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6454) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6769) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24002) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6646) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30837) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27503) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17009) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2922) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14445) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3480) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30351) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6804) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6274) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15393) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13609) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15527) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15922) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5904) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13013) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18259) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17830) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21293) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27247) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8549) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26646) * $signed(input_fmap_85[7:0]) +
	( 14'sd 8042) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22448) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16640) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3391) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30418) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28089) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3218) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32671) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9650) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26849) * $signed(input_fmap_96[7:0]) +
	( 11'sd 554) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20634) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1082) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13608) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14770) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27170) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_106[7:0]) +
	( 11'sd 555) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5196) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19007) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28713) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9003) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8506) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5348) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18794) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6384) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18208) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22324) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5431) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6860) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24492) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9068) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1079) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 15'sd 12087) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25337) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19211) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7753) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15942) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11006) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22620) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9130) * $signed(input_fmap_16[7:0]) +
	( 11'sd 688) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26732) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27751) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24093) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7885) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30601) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2400) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16430) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_30[7:0]) +
	( 10'sd 465) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24536) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4461) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23367) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27987) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4337) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7314) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19701) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21245) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27700) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24593) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5961) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7118) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17322) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22387) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30963) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9261) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15965) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2633) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22083) * $signed(input_fmap_64[7:0]) +
	( 10'sd 447) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25362) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21588) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2542) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31829) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14471) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4849) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8603) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11055) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29751) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25121) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10876) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2146) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32593) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13892) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23579) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10182) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17380) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11814) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26164) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19981) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3490) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9705) * $signed(input_fmap_91[7:0]) +
	( 12'sd 2010) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29885) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20076) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29170) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26177) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28123) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7716) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2149) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2702) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17921) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6976) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7085) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16258) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30954) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17167) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19473) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7840) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3674) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9010) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12300) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17321) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20575) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1571) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12728) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23866) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 12'sd 1687) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_1[7:0]) +
	( 11'sd 823) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16788) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27353) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30145) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6536) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16963) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21337) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26603) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12883) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15637) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31956) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7767) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32017) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3344) * $signed(input_fmap_22[7:0]) +
	( 11'sd 724) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21619) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21789) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17411) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29929) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31313) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4679) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31145) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11220) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23990) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9639) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25839) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31646) * $signed(input_fmap_43[7:0]) +
	( 8'sd 69) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26909) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25860) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22658) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20995) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25618) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27555) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30147) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8859) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15052) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15674) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8745) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20158) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22550) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16426) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10301) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29558) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4325) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16512) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12076) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29370) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15634) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26503) * $signed(input_fmap_80[7:0]) +
	( 11'sd 1007) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1302) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24108) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17561) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22093) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15443) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4732) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1444) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29526) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9241) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23176) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7918) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16821) * $signed(input_fmap_97[7:0]) +
	( 11'sd 708) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23343) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19220) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13115) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16754) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26537) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1939) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21814) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17052) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24388) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29322) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20528) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26824) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20570) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12705) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21159) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5843) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 15'sd 10722) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25959) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17915) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17518) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26546) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20106) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3381) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22566) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18715) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9451) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9334) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13335) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9249) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25316) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4482) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_20[7:0]) +
	( 11'sd 829) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3585) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19581) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9498) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14592) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31595) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_32[7:0]) +
	( 10'sd 457) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10447) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21597) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20793) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16839) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9111) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22521) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17653) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22295) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20788) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16734) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16938) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15867) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7255) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26943) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2312) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18281) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31967) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21681) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1404) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9657) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25648) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9346) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22974) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14099) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12240) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29965) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16106) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28038) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26870) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25921) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13722) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32121) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13108) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16817) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2682) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29379) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14858) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13546) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21502) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29500) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31902) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23748) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2312) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15537) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32327) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22053) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3297) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10066) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28321) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31537) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 12'sd 1584) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3824) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28118) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7276) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12220) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16980) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1332) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22092) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23888) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19986) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6444) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21115) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26504) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10024) * $signed(input_fmap_14[7:0]) +
	( 7'sd 58) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24662) * $signed(input_fmap_16[7:0]) +
	( 9'sd 183) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22469) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7145) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28084) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26356) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9815) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11139) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26920) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22669) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12366) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24528) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14297) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20499) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29620) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31532) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29469) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25012) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10688) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22544) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15652) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19837) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15318) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24433) * $signed(input_fmap_52[7:0]) +
	( 9'sd 174) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25153) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18790) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12057) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9447) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31365) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16921) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23156) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31505) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8642) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30047) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14286) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23703) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24307) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18898) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31233) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4665) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18361) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_80[7:0]) +
	( 9'sd 233) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8779) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_85[7:0]) +
	( 11'sd 605) * $signed(input_fmap_86[7:0]) +
	( 9'sd 177) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16781) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15466) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24856) * $signed(input_fmap_91[7:0]) +
	( 7'sd 44) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30195) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1507) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26324) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8489) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27050) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4665) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9827) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11396) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23351) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6743) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3702) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_111[7:0]) +
	( 11'sd 647) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5103) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12493) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16725) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15513) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11301) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10394) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3962) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28378) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9221) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6649) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16460) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10968) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1178) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 16'sd 29038) * $signed(input_fmap_0[7:0]) +
	( 14'sd 8033) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3492) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6968) * $signed(input_fmap_3[7:0]) +
	( 13'sd 4082) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16857) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6599) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3431) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24584) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5401) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5273) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4561) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4453) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21364) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30451) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3912) * $signed(input_fmap_20[7:0]) +
	( 9'sd 167) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26253) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11653) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29248) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19115) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7753) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28571) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30551) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30964) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10240) * $signed(input_fmap_36[7:0]) +
	( 7'sd 46) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1429) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2402) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28517) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30474) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14599) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11925) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25387) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4765) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9618) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7660) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11773) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6343) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28403) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15143) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_59[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27061) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27663) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15165) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14127) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2749) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13371) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7253) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14287) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22104) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26367) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12566) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8774) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9918) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15710) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2052) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5621) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9528) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3934) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10472) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1071) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2051) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3430) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12530) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16494) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3195) * $signed(input_fmap_98[7:0]) +
	( 11'sd 997) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5492) * $signed(input_fmap_100[7:0]) +
	( 9'sd 241) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18607) * $signed(input_fmap_102[7:0]) +
	( 11'sd 600) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27882) * $signed(input_fmap_106[7:0]) +
	( 10'sd 449) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31653) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6131) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23295) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7096) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11677) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29598) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3874) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26579) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_123[7:0]) +
	( 10'sd 378) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18597) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12254) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 15'sd 9010) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31247) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24942) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14453) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29756) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14084) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25284) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20100) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11781) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27528) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21929) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23720) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23584) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8477) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24922) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2709) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29640) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31686) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9014) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14106) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23449) * $signed(input_fmap_31[7:0]) +
	( 10'sd 353) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28682) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18023) * $signed(input_fmap_35[7:0]) +
	( 9'sd 145) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9693) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1780) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6229) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4326) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21976) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6686) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16234) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1970) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25560) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6068) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8570) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_54[7:0]) +
	( 10'sd 495) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29442) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15539) * $signed(input_fmap_58[7:0]) +
	( 11'sd 586) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11748) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4727) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19999) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1284) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4676) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31139) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6386) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14858) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17903) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24893) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4488) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24948) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32293) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15299) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30678) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10548) * $signed(input_fmap_90[7:0]) +
	( 9'sd 190) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30004) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19147) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15137) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18570) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2167) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_97[7:0]) +
	( 13'sd 4028) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28505) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10250) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3979) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3677) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27136) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13697) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25102) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3288) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14980) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20323) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5435) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28264) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28254) * $signed(input_fmap_116[7:0]) +
	( 12'sd 2036) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5360) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11665) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21950) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5358) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25830) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8248) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23156) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 16'sd 27820) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18878) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27844) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1187) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25091) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31551) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23336) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1411) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11093) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4611) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31694) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8120) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_20[7:0]) +
	( 11'sd 598) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31365) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2847) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5216) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17477) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27393) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13227) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18430) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7746) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_35[7:0]) +
	( 11'sd 898) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28829) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2212) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11413) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28380) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31323) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6540) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29454) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18995) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24749) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19450) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5710) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29187) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28579) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18600) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25881) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28595) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20857) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11720) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13267) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31893) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10039) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19104) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10542) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10157) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30976) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1202) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31349) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12062) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18732) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27014) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8453) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7327) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16398) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18696) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30193) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30710) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8030) * $signed(input_fmap_88[7:0]) +
	( 11'sd 753) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11050) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19744) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23923) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13645) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4589) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23493) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12317) * $signed(input_fmap_98[7:0]) +
	( 10'sd 372) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29252) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19517) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16476) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16593) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3926) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31096) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7352) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13520) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26414) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28691) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24619) * $signed(input_fmap_118[7:0]) +
	( 11'sd 698) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14451) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14367) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2202) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27276) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 16'sd 20468) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3077) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32231) * $signed(input_fmap_2[7:0]) +
	( 9'sd 220) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5452) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30567) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23600) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24077) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28508) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22291) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28513) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22149) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_19[7:0]) +
	( 7'sd 36) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8101) * $signed(input_fmap_27[7:0]) +
	( 9'sd 203) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9071) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20189) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19818) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5508) * $signed(input_fmap_32[7:0]) +
	( 11'sd 689) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19925) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20668) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29557) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21318) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24481) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4717) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16008) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32496) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5173) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5309) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19328) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27183) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3040) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6475) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1416) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3435) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27826) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19644) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16963) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11268) * $signed(input_fmap_61[7:0]) +
	( 11'sd 544) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21088) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20481) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30933) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1106) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25711) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8319) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14486) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3574) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19400) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12291) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5907) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6599) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29088) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29226) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4267) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30585) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31906) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30151) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9888) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30202) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13070) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5243) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27802) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6085) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20436) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29335) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17030) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28762) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25054) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31839) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23526) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19242) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31649) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26219) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12022) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_119[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17546) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6802) * $signed(input_fmap_123[7:0]) +
	( 9'sd 154) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18731) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31253) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9937) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 16'sd 32159) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19837) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21874) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32578) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1319) * $signed(input_fmap_7[7:0]) +
	( 11'sd 981) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25604) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14845) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17032) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_12[7:0]) +
	( 10'sd 470) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3741) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21652) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16075) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20819) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5058) * $signed(input_fmap_21[7:0]) +
	( 9'sd 148) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14833) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22721) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3801) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27685) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22001) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29286) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16960) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18343) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20204) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29457) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32515) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27930) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17788) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26097) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4568) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25722) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1043) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10956) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16565) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2544) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8291) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3843) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11320) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18923) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20327) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23518) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2211) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22032) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31928) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10698) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13954) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28075) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27699) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4370) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12163) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19755) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12835) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27562) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9983) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1885) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13923) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25033) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2337) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20834) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8914) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1903) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24711) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10745) * $signed(input_fmap_99[7:0]) +
	( 10'sd 416) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10641) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6270) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23662) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23710) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30728) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26508) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6796) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1476) * $signed(input_fmap_114[7:0]) +
	( 11'sd 652) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6351) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25324) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17043) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30622) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10940) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9961) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27126) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8530) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31189) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 15'sd 13402) * $signed(input_fmap_0[7:0]) +
	( 10'sd 504) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19449) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1543) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14398) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13828) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27803) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28251) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6461) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18150) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1770) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31955) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29316) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4777) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29096) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1752) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17712) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29929) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15435) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_28[7:0]) +
	( 11'sd 582) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4205) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6264) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10645) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21933) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26798) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_37[7:0]) +
	( 11'sd 866) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7509) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10943) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17035) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27551) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25767) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10610) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2930) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5732) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6770) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6285) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_57[7:0]) +
	( 9'sd 249) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16038) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31685) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2176) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12598) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24481) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29346) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29054) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30189) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29306) * $signed(input_fmap_68[7:0]) +
	( 11'sd 725) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16547) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8819) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21112) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4597) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13761) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1527) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11531) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13437) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31794) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11826) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3290) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5207) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17256) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11105) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4377) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24021) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22741) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19774) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15568) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15028) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23910) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18457) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30655) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31707) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17506) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28235) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5781) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15374) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22840) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5635) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27412) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29504) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26027) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29071) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15343) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19572) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12568) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20441) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2097) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11165) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9005) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4973) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 16'sd 30769) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21064) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18641) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17642) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7866) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2171) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15611) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20602) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10418) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13804) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7889) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26791) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29593) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26440) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15930) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22511) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8563) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12104) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4567) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2520) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2362) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26436) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30765) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7746) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5451) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20558) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14251) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5394) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16877) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5450) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28192) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10639) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11022) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_53[7:0]) +
	( 8'sd 77) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22824) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12935) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10560) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27182) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1644) * $signed(input_fmap_62[7:0]) +
	( 11'sd 1022) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_65[7:0]) +
	( 11'sd 568) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15764) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25400) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23600) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21976) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17101) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25550) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14242) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11330) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21336) * $signed(input_fmap_80[7:0]) +
	( 11'sd 861) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23392) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31847) * $signed(input_fmap_84[7:0]) +
	( 11'sd 564) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26752) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27683) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15045) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22931) * $signed(input_fmap_91[7:0]) +
	( 10'sd 446) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16854) * $signed(input_fmap_93[7:0]) +
	( 6'sd 26) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30822) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24577) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15750) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30167) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30023) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6933) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1406) * $signed(input_fmap_106[7:0]) +
	( 11'sd 853) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21085) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26646) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13597) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24147) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26788) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9389) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23158) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1345) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28988) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20789) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14928) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13640) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 16'sd 23157) * $signed(input_fmap_0[7:0]) +
	( 10'sd 405) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14726) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2240) * $signed(input_fmap_3[7:0]) +
	( 11'sd 547) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_5[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2580) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10311) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1584) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25033) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11251) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8877) * $signed(input_fmap_16[7:0]) +
	( 11'sd 709) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7857) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29833) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20707) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11999) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13337) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21988) * $signed(input_fmap_24[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8581) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7023) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8183) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5617) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28559) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29295) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9677) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19826) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16956) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10994) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13546) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25237) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24561) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10104) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15015) * $signed(input_fmap_55[7:0]) +
	( 13'sd 4010) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32687) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28903) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1325) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14698) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17391) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9794) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5152) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7409) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15635) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28470) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31386) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31537) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15852) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19497) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6967) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3917) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26701) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11818) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5717) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2944) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17578) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13393) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25555) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5504) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3941) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30271) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25861) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18419) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28165) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3726) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1107) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20929) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26073) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31068) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15247) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 15'sd 9076) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26340) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20100) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29314) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28172) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30726) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22259) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29761) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18454) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2734) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18829) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5031) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28507) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22161) * $signed(input_fmap_25[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5807) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23370) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17327) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9733) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29119) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14346) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18894) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10095) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12673) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13664) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30798) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9982) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19892) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24208) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20664) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12627) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7044) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22652) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26777) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14765) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7125) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3154) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29673) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14864) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26019) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3768) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29052) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3252) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9906) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29733) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9405) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13730) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12967) * $signed(input_fmap_74[7:0]) +
	( 14'sd 8084) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20707) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13055) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32102) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29045) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_82[7:0]) +
	( 14'sd 8160) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1575) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4926) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14540) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5395) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16486) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17387) * $signed(input_fmap_102[7:0]) +
	( 10'sd 295) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24629) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21537) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8080) * $signed(input_fmap_111[7:0]) +
	( 9'sd 136) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9947) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29768) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3110) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13433) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10480) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26303) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19791) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26057) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24354) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22923) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1037) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 16'sd 30406) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27703) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27636) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17769) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29501) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18084) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12810) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4232) * $signed(input_fmap_12[7:0]) +
	( 9'sd 169) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_15[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4772) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1555) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29837) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22372) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30952) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30506) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2293) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6154) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3308) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26601) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32012) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_31[7:0]) +
	( 10'sd 491) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18826) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27471) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15865) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8836) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6199) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17239) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_45[7:0]) +
	( 10'sd 262) * $signed(input_fmap_46[7:0]) +
	( 11'sd 576) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26950) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15559) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7924) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18286) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6043) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26519) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5038) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21040) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9889) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1751) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26632) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31319) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24725) * $signed(input_fmap_67[7:0]) +
	( 9'sd 161) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1106) * $signed(input_fmap_69[7:0]) +
	( 9'sd 248) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2703) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20649) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18167) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22763) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25093) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4504) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26619) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4997) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1390) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13621) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13924) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_94[7:0]) +
	( 8'sd 85) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26164) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25890) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22721) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17936) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13967) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9819) * $signed(input_fmap_107[7:0]) +
	( 11'sd 611) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27794) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16690) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23594) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14377) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24122) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5442) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25187) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20683) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31275) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7737) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25974) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23411) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12656) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7545) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3827) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 15'sd 10134) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14804) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20245) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17460) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5991) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9995) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11597) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31759) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6052) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15949) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29340) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14632) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26729) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21364) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9469) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2981) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17893) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21045) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7370) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11727) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14467) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9358) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29144) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12763) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10563) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12617) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18003) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32725) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23749) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9517) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30050) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3136) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7675) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22542) * $signed(input_fmap_51[7:0]) +
	( 12'sd 2013) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28064) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21811) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26435) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3451) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3626) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24243) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10433) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23832) * $signed(input_fmap_65[7:0]) +
	( 13'sd 4027) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10346) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30451) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7542) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24389) * $signed(input_fmap_71[7:0]) +
	( 14'sd 8104) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28973) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1287) * $signed(input_fmap_76[7:0]) +
	( 12'sd 2004) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11797) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7904) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21705) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6172) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3643) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2202) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7830) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25940) * $signed(input_fmap_86[7:0]) +
	( 4'sd 4) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21066) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26196) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12990) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10318) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17820) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24606) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27626) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5441) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5573) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31604) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18372) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15843) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9633) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25284) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20239) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13380) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22183) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3488) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10529) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13932) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8730) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3904) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28559) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4694) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22324) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12795) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26259) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21846) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1706) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 10'sd 405) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13912) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12331) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23645) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2925) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9552) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16986) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27290) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26805) * $signed(input_fmap_12[7:0]) +
	( 14'sd 8095) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17528) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13915) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29920) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29418) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28654) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16257) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14475) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24638) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9698) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14778) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22195) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6790) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20086) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26068) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23650) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17501) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31157) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1026) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29913) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27651) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13518) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16736) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8361) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25294) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4784) * $signed(input_fmap_44[7:0]) +
	( 10'sd 464) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31187) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1169) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7038) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28069) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17103) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18161) * $signed(input_fmap_52[7:0]) +
	( 13'sd 4081) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27903) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3166) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4716) * $signed(input_fmap_58[7:0]) +
	( 10'sd 277) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20861) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7341) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28599) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1341) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29462) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8573) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31549) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20108) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2920) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23887) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18126) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8946) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25226) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15281) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10151) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3524) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7177) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11425) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22279) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11536) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1497) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20463) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6891) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9821) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17789) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26442) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27012) * $signed(input_fmap_105[7:0]) +
	( 11'sd 656) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30845) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17410) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5325) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22580) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17424) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29884) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25844) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24492) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28378) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7611) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1416) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4895) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15922) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26159) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23777) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2093) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 16'sd 29979) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14906) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9582) * $signed(input_fmap_6[7:0]) +
	( 11'sd 959) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15839) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15188) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12579) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1066) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31797) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11988) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8817) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1958) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21960) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22046) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32252) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18491) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7783) * $signed(input_fmap_32[7:0]) +
	( 9'sd 221) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10031) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31590) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10892) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12503) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15565) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25667) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18723) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15852) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10092) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30361) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14817) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29979) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7821) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23308) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28612) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29840) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22816) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5712) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21635) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11823) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30891) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7285) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4618) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_70[7:0]) +
	( 10'sd 360) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17742) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21067) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24113) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21244) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10218) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20533) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5058) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21632) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22387) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22768) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_86[7:0]) +
	( 10'sd 495) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29699) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5019) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7711) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10156) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21933) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15147) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19086) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4129) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10995) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6907) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28961) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15185) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19137) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7320) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24951) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29205) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9834) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30581) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8788) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27562) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1958) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17378) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23352) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 14'sd 7290) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25076) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16435) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2160) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9591) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26560) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15003) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26726) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22145) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1654) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24879) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27445) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9133) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21913) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1669) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2182) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4829) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25335) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10619) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29353) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24480) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25580) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11845) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8393) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12613) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11010) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29371) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22824) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14804) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26708) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28243) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26796) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21341) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1821) * $signed(input_fmap_47[7:0]) +
	( 11'sd 555) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14478) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14790) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15276) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8893) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31073) * $signed(input_fmap_56[7:0]) +
	( 11'sd 929) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16035) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11240) * $signed(input_fmap_60[7:0]) +
	( 10'sd 388) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6841) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11169) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31988) * $signed(input_fmap_66[7:0]) +
	( 10'sd 292) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7477) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12852) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28533) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32074) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1148) * $signed(input_fmap_75[7:0]) +
	( 11'sd 585) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7185) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7339) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27889) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19360) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11037) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17981) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9521) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22617) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11263) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6581) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25667) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8181) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1826) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27169) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7528) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32386) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28286) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28860) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30590) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24623) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10486) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20093) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9934) * $signed(input_fmap_103[7:0]) +
	( 8'sd 84) * $signed(input_fmap_104[7:0]) +
	( 10'sd 486) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25300) * $signed(input_fmap_106[7:0]) +
	( 12'sd 2002) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4838) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7284) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3397) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32336) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19745) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12171) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21783) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7693) * $signed(input_fmap_120[7:0]) +
	( 7'sd 63) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10529) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12511) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1376) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26870) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 15'sd 16174) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12062) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24274) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30934) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21083) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19407) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18186) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26346) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25076) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8788) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10670) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2502) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20745) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18383) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18837) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8605) * $signed(input_fmap_20[7:0]) +
	( 11'sd 575) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32209) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12822) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15371) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32062) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30155) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22008) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26974) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7534) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_37[7:0]) +
	( 11'sd 714) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16546) * $signed(input_fmap_42[7:0]) +
	( 11'sd 624) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5308) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29568) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9767) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31461) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25474) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29372) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1926) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6061) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25071) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22150) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3752) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15580) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10125) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13899) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25023) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25328) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9505) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21420) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13948) * $signed(input_fmap_71[7:0]) +
	( 10'sd 326) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6111) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6703) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25461) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30592) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4224) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14338) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2805) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10387) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30153) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27318) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18224) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32231) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27697) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14309) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18416) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14738) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32097) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30194) * $signed(input_fmap_102[7:0]) +
	( 10'sd 385) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28484) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20360) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5250) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2789) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7595) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4729) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11550) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29019) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23944) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28141) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5883) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10565) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30848) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21994) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9236) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22344) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 14'sd 4196) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3641) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22120) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_4[7:0]) +
	( 11'sd 773) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26366) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_7[7:0]) +
	( 10'sd 270) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5185) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5263) * $signed(input_fmap_13[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28999) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6112) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26516) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_20[7:0]) +
	( 9'sd 209) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14879) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16051) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6059) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_27[7:0]) +
	( 11'sd 786) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12586) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3371) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27762) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17866) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25097) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20782) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12996) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7681) * $signed(input_fmap_40[7:0]) +
	( 11'sd 798) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8168) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26158) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8278) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6081) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12650) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18976) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19002) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14918) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25061) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18846) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5527) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8205) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27174) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19215) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25374) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12165) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18101) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8677) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24407) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15206) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19145) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3379) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22205) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28269) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14530) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16276) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20361) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1905) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12463) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22537) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21358) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27494) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5530) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29542) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7864) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16151) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29267) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9986) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6151) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16111) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12330) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_120[7:0]) +
	( 7'sd 54) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8903) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16768) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 15'sd 8369) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23016) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8771) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11258) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26507) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10637) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3620) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12819) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16814) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31149) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10387) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26769) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3444) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13553) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10736) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5005) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22691) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1306) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26893) * $signed(input_fmap_34[7:0]) +
	( 11'sd 886) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1570) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30336) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1306) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15496) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28618) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8404) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24245) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13485) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27646) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26596) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3767) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18173) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26029) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12578) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15956) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26281) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4297) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2184) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8543) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27132) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18275) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24158) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29058) * $signed(input_fmap_72[7:0]) +
	( 11'sd 649) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20553) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12039) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28747) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2332) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6929) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14146) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3486) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6934) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22363) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4759) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21215) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20442) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7823) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2921) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9864) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11109) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6664) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15262) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31654) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22142) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20882) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16708) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23339) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9513) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_110[7:0]) +
	( 8'sd 104) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28067) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11714) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31561) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25814) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24511) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15525) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26873) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13107) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9887) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19929) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25577) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8330) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 15'sd 9245) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21713) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18923) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10410) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15002) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16349) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22207) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13579) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26917) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26197) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30149) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2677) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26016) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16689) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16224) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25779) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20000) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28715) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15350) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28690) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25261) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31244) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20500) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21300) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15919) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27857) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6106) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7389) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12607) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15921) * $signed(input_fmap_46[7:0]) +
	( 7'sd 60) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20986) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13423) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_51[7:0]) +
	( 9'sd 131) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9983) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5193) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15561) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4510) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5132) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10529) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14505) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30410) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4407) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23973) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4431) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6896) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12283) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15308) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13524) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29332) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31558) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4681) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31222) * $signed(input_fmap_84[7:0]) +
	( 11'sd 960) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20268) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24830) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13165) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24477) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30929) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15591) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19979) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31011) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21617) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24720) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21353) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31149) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31876) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1155) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31480) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23870) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32460) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28161) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14196) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12595) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6755) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11009) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1946) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7132) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25735) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30104) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25519) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_120[7:0]) +
	( 10'sd 359) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30336) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11229) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24337) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 16'sd 29492) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27845) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7068) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28390) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2375) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5871) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14948) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17475) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30348) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28125) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14345) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26279) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21293) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1915) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11724) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29043) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28611) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26092) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19778) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1798) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29495) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16219) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9108) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15727) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3181) * $signed(input_fmap_36[7:0]) +
	( 9'sd 178) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7542) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15897) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28116) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11394) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15944) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15261) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15463) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26376) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22639) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6392) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11522) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17043) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4242) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29812) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16183) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22689) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3523) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21192) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30057) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18778) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16357) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6621) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31500) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30215) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32573) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14279) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4547) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1798) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25485) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23079) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25253) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24836) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7279) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16780) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23460) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18341) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16991) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10470) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10355) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23761) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22424) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23513) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14093) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11196) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4306) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17184) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26231) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17741) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26867) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5336) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3371) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21388) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2723) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4687) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18244) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28928) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30021) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 16'sd 32711) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6476) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31258) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6355) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5232) * $signed(input_fmap_5[7:0]) +
	( 11'sd 590) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19817) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31283) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21324) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2996) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26777) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14659) * $signed(input_fmap_20[7:0]) +
	( 13'sd 4004) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30662) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14160) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7722) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4242) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13988) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23691) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18832) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16955) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31972) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6414) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21424) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3860) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31995) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16877) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3336) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3167) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1343) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3507) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6308) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11715) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18818) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17572) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9026) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32464) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31919) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11984) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1707) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14525) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1521) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16991) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5978) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7582) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19132) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9312) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1116) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25795) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22354) * $signed(input_fmap_74[7:0]) +
	( 11'sd 684) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2933) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26553) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25032) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29568) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16744) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20094) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1040) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6253) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2910) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2469) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9124) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28466) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26121) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16396) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32054) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26947) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25798) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11447) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22035) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_102[7:0]) +
	( 8'sd 88) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22783) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26372) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22419) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10546) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29899) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16418) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17818) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6139) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24739) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26536) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6750) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23633) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30155) * $signed(input_fmap_124[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 16'sd 26219) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8381) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22512) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6364) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9268) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6268) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10317) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25032) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12841) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1358) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10417) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20868) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9894) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13422) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25391) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26525) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3330) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3234) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_23[7:0]) +
	( 10'sd 357) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10341) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16473) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21471) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7115) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27051) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28268) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13668) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13108) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11435) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5553) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28993) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_42[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11994) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27184) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12331) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13750) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5633) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25287) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4747) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8618) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12530) * $signed(input_fmap_54[7:0]) +
	( 9'sd 211) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26884) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3607) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30476) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21255) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20516) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8762) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7385) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15174) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16152) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29923) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23559) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7722) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8357) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30979) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4476) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2848) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5142) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10242) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31443) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8276) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7698) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7391) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26793) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29507) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8773) * $signed(input_fmap_90[7:0]) +
	( 11'sd 1021) * $signed(input_fmap_91[7:0]) +
	( 9'sd 153) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19744) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2592) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30907) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22218) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6000) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10212) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4871) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30725) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1476) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31401) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22228) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7501) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31983) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32295) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6899) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4559) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18613) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17096) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30776) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5988) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20328) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16662) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24676) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 16'sd 21729) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30710) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27331) * $signed(input_fmap_2[7:0]) +
	( 11'sd 604) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30688) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29041) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21757) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16533) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29814) * $signed(input_fmap_8[7:0]) +
	( 11'sd 710) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11495) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30184) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14099) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25006) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10647) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1204) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11640) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31173) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10202) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18453) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10437) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10365) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28035) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21287) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15019) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4521) * $signed(input_fmap_34[7:0]) +
	( 5'sd 9) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8556) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1484) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22504) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23699) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12199) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23467) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14604) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25224) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13906) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18276) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10033) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22579) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13996) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20727) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14146) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27823) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28346) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23018) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28774) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29516) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28858) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9552) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_75[7:0]) +
	( 11'sd 543) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31057) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16691) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14836) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5010) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26662) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1626) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4337) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1904) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4195) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11275) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32632) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11788) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26442) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20518) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19254) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19222) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29241) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29274) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22922) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20836) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25208) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16957) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10313) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26413) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22420) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2346) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24992) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19949) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5942) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26962) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27246) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 14'sd 7682) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8282) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32226) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13977) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30895) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12857) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32067) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1358) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5670) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24637) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23124) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18701) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27388) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26261) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21631) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28023) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26738) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16730) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5833) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12439) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9846) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19431) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10200) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26144) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7313) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14248) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3316) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13495) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5009) * $signed(input_fmap_41[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27074) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30642) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11151) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13139) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10223) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29780) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18358) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7771) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30678) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9962) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18168) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26673) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6934) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20261) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4171) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32187) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18815) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24515) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25647) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14495) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29960) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1989) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25885) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1926) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23574) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24843) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23708) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_87[7:0]) +
	( 10'sd 459) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6524) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25148) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31043) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23084) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7681) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24348) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9349) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_98[7:0]) +
	( 11'sd 818) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4742) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14080) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19081) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28516) * $signed(input_fmap_103[7:0]) +
	( 11'sd 941) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1730) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9719) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32593) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20193) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26254) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16561) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30757) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17406) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3112) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16595) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26392) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 13'sd 2983) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19611) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21860) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2315) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23848) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2334) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1232) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21269) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4762) * $signed(input_fmap_11[7:0]) +
	( 14'sd 8130) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15203) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5074) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19399) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1441) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3248) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5363) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4514) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24380) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7115) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21080) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_23[7:0]) +
	( 14'sd 8040) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2778) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26326) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23882) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12779) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3370) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21831) * $signed(input_fmap_31[7:0]) +
	( 5'sd 14) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22510) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1312) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21157) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3528) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5302) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13622) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11603) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19523) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21355) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12313) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3754) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7159) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7919) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21415) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18395) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8224) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17766) * $signed(input_fmap_57[7:0]) +
	( 8'sd 95) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32245) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16573) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19259) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12540) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32084) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22211) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12721) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10648) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12503) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9273) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5547) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6244) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25676) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10298) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2960) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2904) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14988) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28047) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13900) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16045) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1229) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2348) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13616) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_91[7:0]) +
	( 11'sd 694) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29639) * $signed(input_fmap_94[7:0]) +
	( 11'sd 997) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32074) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13933) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5219) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11197) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2142) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14823) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27578) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10706) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14865) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15484) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18412) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4492) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30108) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11358) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30682) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13486) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2147) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15129) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 15'sd 10245) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13358) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28093) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22160) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2566) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8386) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11443) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20797) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31191) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2052) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1397) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7944) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9441) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5308) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23749) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15687) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17809) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18572) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27408) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28675) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19860) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21316) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15394) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8495) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2254) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17764) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17231) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4740) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5585) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1148) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_46[7:0]) +
	( 11'sd 852) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4916) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1690) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9377) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14159) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23066) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31230) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10241) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7943) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27552) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23596) * $signed(input_fmap_61[7:0]) +
	( 10'sd 310) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14321) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9056) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11096) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13859) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2572) * $signed(input_fmap_68[7:0]) +
	( 11'sd 877) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12555) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2703) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30513) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6450) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12675) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25362) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31266) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14747) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4542) * $signed(input_fmap_87[7:0]) +
	( 9'sd 133) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28901) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7429) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13334) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23400) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28758) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32184) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16363) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22071) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4893) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21319) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11562) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3944) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9616) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25331) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11844) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4608) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2878) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9601) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17472) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1203) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1858) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29065) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17252) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5773) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 14'sd 4167) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3199) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3391) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18178) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5545) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8388) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7246) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32068) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19522) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15176) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1175) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20369) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3351) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27146) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19895) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5936) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10712) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18101) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17286) * $signed(input_fmap_23[7:0]) +
	( 7'sd 36) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4539) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25776) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17862) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28534) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27013) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22689) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10877) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1326) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16759) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6328) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22778) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4516) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13084) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14535) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25202) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13726) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17353) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31176) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24967) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5244) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30296) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21452) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20575) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14868) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18274) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30076) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18029) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32211) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7839) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31093) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10534) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21291) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1761) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20341) * $signed(input_fmap_78[7:0]) +
	( 10'sd 503) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14299) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16354) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10636) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16264) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15245) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10993) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19979) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6124) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12601) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27507) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23180) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24452) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30082) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21975) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16386) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17994) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13168) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3746) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15355) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20834) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14340) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7349) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3230) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2211) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6578) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13296) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14956) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 15'sd 13866) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31995) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22131) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31691) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19530) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2195) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18662) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5320) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8400) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23163) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16898) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21310) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19536) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17373) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10403) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26841) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32562) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11709) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18719) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21021) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18569) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12172) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17330) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18184) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21642) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14092) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16098) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4639) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3936) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9083) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20398) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11326) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13138) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26059) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32114) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21918) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9847) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22584) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26175) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16582) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20998) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14037) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10781) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13837) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14106) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29273) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29208) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18453) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18945) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29999) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30757) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12589) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1145) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19505) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5329) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9210) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13055) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29035) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17704) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28335) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23002) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32365) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27704) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20145) * $signed(input_fmap_94[7:0]) +
	( 11'sd 674) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2657) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_99[7:0]) +
	( 11'sd 787) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3098) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7827) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7386) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6675) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15655) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5207) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24357) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9644) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21367) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19183) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22749) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7904) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1109) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22602) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28704) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 16'sd 27998) * $signed(input_fmap_0[7:0]) +
	( 11'sd 562) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12842) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30943) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3291) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13459) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32201) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22969) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26722) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16432) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26932) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15079) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27057) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4605) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27246) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8283) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4528) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5465) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29989) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27226) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18468) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22465) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12395) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25205) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27305) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19080) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25764) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4684) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23886) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3296) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10398) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17923) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3546) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18752) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11948) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32551) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27589) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_62[7:0]) +
	( 10'sd 433) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7884) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9433) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2406) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10919) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15499) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17086) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16872) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9795) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6509) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32521) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9504) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24208) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19330) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3088) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3729) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24483) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17248) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25502) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22709) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26018) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21725) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9873) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24908) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13740) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12305) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29511) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11834) * $signed(input_fmap_110[7:0]) +
	( 10'sd 446) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13061) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11427) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4668) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13344) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17315) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22751) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15138) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17682) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16384) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29256) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11304) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21513) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19002) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9139) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 14'sd 7310) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22395) * $signed(input_fmap_1[7:0]) +
	( 11'sd 573) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22137) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13692) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32409) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_9[7:0]) +
	( 10'sd 375) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19600) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19150) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13562) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1842) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22718) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17616) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19289) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1937) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11935) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17198) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6169) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24730) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20386) * $signed(input_fmap_29[7:0]) +
	( 11'sd 986) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10845) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24261) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31283) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29609) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30150) * $signed(input_fmap_37[7:0]) +
	( 11'sd 830) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21152) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14048) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1560) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5855) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15388) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31196) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1535) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22193) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12471) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10699) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22566) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22378) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3266) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24262) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27737) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12536) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14460) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10348) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3947) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6413) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8581) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12949) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1345) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15121) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22572) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6450) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18035) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31713) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30042) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29148) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26265) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31448) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8859) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2747) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25196) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27153) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29192) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14956) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4430) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19799) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21302) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26410) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21696) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4441) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23976) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3606) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2934) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31620) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15886) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 14'sd 8093) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1465) * $signed(input_fmap_1[7:0]) +
	( 11'sd 714) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14305) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10387) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1560) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31324) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13053) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22472) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6032) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5651) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17379) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6362) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16880) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26117) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29887) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5496) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22228) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32057) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7473) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20068) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3565) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18277) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22518) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8274) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23279) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1259) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26086) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20756) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29848) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16845) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3659) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7879) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31650) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5083) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26426) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6449) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20911) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2090) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32538) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12794) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18903) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23147) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26332) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9908) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27600) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12349) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13640) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27224) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14427) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31256) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18805) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26692) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19974) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31063) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7979) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11069) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19431) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9779) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5710) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27687) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16079) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10418) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27353) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19214) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5637) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3315) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1686) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28906) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32289) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14457) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3128) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7462) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25290) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11753) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1633) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5604) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17640) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30695) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19119) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 15'sd 8897) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5855) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19360) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30254) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1774) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21096) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12390) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16586) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28499) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1775) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27703) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20028) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17725) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12201) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4324) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5595) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12712) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21478) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4487) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29047) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7200) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25029) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1132) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2752) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22270) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16722) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15695) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22002) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10232) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20609) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17815) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13109) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23003) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30687) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28115) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5517) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31099) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17251) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2747) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32161) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11648) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23037) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30614) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26922) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15759) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29630) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27992) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31277) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14551) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28878) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27657) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30612) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9049) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25544) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19929) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2984) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1530) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6717) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7727) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5298) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25801) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2105) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22688) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9027) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15769) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32175) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8824) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3763) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24970) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11884) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23186) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22096) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24708) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12746) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32177) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29407) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31361) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8472) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13049) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23895) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7496) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26701) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18030) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6108) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_124[7:0]) +
	( 11'sd 995) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24480) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 16'sd 25459) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6530) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7029) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24429) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4880) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11657) * $signed(input_fmap_9[7:0]) +
	( 8'sd 126) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4823) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16928) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15698) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32719) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23968) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15947) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10227) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4717) * $signed(input_fmap_19[7:0]) +
	( 11'sd 814) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20111) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13228) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23639) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29121) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30558) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_32[7:0]) +
	( 10'sd 447) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4442) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25015) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23334) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17543) * $signed(input_fmap_39[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31629) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29417) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23777) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31530) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11798) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15653) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4492) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17813) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14947) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9423) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16834) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30380) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18224) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28578) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32096) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31582) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26903) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21189) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22995) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28714) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21573) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4325) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28945) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30621) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17032) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11850) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22604) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13927) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5282) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10527) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15336) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1416) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1112) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30954) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25846) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17647) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23159) * $signed(input_fmap_95[7:0]) +
	( 11'sd 583) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16532) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7019) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14311) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6904) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19379) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15410) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11361) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18519) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7382) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14957) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13903) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6576) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8489) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23241) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23326) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6217) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26580) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8179) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 15'sd 11919) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15655) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7434) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16263) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1231) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9019) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23413) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15095) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31341) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2798) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21548) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9584) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24297) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8232) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23238) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2390) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19127) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14572) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22679) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7215) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_36[7:0]) +
	( 13'sd 4070) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29424) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28846) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15666) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24641) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19337) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23308) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28175) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8653) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14911) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23848) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32562) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21586) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9798) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21834) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12621) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3319) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32590) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24110) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15281) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2859) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26351) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18911) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7207) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13358) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11998) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10894) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5560) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17506) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25252) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_81[7:0]) +
	( 10'sd 256) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15218) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14108) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22530) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24962) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16140) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28198) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5943) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1855) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8133) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18807) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20922) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25734) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31122) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30385) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25088) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8794) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20219) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19638) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5247) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28583) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9585) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7915) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24573) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24142) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14654) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13590) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6591) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32502) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 16'sd 21530) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1280) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11388) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20951) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20733) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13738) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8833) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13583) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11071) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15580) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26720) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19337) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2871) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29655) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2890) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30409) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1131) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25101) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18188) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31878) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23936) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19535) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1740) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21822) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27347) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3099) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21279) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16414) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20570) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14300) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10782) * $signed(input_fmap_45[7:0]) +
	( 11'sd 907) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4413) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12900) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14176) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22211) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24689) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12288) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1671) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19109) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11595) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29334) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19924) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10056) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5272) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4270) * $signed(input_fmap_62[7:0]) +
	( 5'sd 8) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21548) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19264) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19259) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9032) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10583) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7033) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19031) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25500) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10100) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16763) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17974) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7119) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25028) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27095) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27099) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29381) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28163) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10083) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_96[7:0]) +
	( 13'sd 4084) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22504) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7948) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11183) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17152) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26866) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16987) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9060) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13017) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6580) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27154) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5538) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2702) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23804) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13861) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23688) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19672) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19035) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 16'sd 30840) * $signed(input_fmap_0[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10734) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6841) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30915) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10865) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1570) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24368) * $signed(input_fmap_10[7:0]) +
	( 11'sd 881) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32124) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17627) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17995) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16192) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4348) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1607) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28979) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25546) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30464) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2890) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26949) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31912) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18392) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8544) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16857) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19283) * $signed(input_fmap_35[7:0]) +
	( 10'sd 378) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19894) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6691) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8655) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25191) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13849) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16580) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19505) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6435) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31547) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27747) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25690) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11973) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11196) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12415) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29617) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18358) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13454) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31900) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19033) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8622) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1593) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32732) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20404) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9329) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18554) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23964) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4398) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12055) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8410) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27071) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23841) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7262) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16640) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28642) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_84[7:0]) +
	( 14'sd 8019) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2876) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22478) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23809) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27724) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31890) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21983) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29891) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23830) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16018) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1055) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17256) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31382) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24538) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11010) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28736) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24599) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21503) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15010) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10298) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25406) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17963) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29699) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13267) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2347) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 15'sd 9608) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22643) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31706) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2392) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32200) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20148) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18533) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7863) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22665) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30139) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3714) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13184) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2808) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10351) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_25[7:0]) +
	( 7'sd 47) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25285) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6854) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15485) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13752) * $signed(input_fmap_31[7:0]) +
	( 11'sd 815) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1671) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26554) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22274) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22992) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25718) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5076) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30168) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31520) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25313) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_46[7:0]) +
	( 10'sd 510) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13837) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22175) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25265) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27412) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28046) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12947) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32011) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15463) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4580) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26635) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32040) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7506) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25755) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26320) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12256) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16512) * $signed(input_fmap_69[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9325) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1605) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7696) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5674) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30536) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4277) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_78[7:0]) +
	( 11'sd 751) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1271) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16672) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26644) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1743) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32071) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11677) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27381) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20794) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22015) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31146) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6024) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1600) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23734) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29412) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30562) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4957) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21585) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23310) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9159) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1142) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30215) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8988) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10223) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19363) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19327) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25305) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21622) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 15'sd 13023) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7525) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23752) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31047) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30560) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27353) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31049) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16913) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26159) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11239) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16340) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28454) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3711) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13465) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9327) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30868) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30657) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32041) * $signed(input_fmap_24[7:0]) +
	( 11'sd 896) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20806) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28687) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32404) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21014) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16744) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10597) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17946) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29367) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25026) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6448) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24824) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24335) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12063) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20419) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20756) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21017) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24376) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15454) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17008) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23017) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6125) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13754) * $signed(input_fmap_60[7:0]) +
	( 10'sd 490) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10005) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29685) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14302) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12336) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31774) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4178) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5120) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30296) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23526) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3683) * $signed(input_fmap_74[7:0]) +
	( 11'sd 899) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21003) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_77[7:0]) +
	( 8'sd 73) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5239) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6954) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24137) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17952) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23549) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11118) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11962) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11407) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29073) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28542) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17115) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2169) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7021) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26653) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8909) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2744) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21746) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24723) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27205) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17452) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23791) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27561) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9843) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6140) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6045) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16434) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21934) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8794) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6043) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21460) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6379) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7838) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27867) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 15'sd 11101) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30925) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28406) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12680) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2882) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31944) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23776) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30936) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12281) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28172) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11316) * $signed(input_fmap_17[7:0]) +
	( 10'sd 303) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14732) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9967) * $signed(input_fmap_22[7:0]) +
	( 11'sd 539) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13242) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5093) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5211) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25910) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19409) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29599) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13746) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29806) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21823) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19303) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13963) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13250) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26848) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8684) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3573) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10355) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11015) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31409) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21961) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15077) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23523) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26453) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4439) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5081) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15860) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21734) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31402) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18457) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21495) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20748) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7781) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17330) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26150) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18813) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21841) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19882) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6291) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18629) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4792) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31795) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12585) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2660) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20632) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1609) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24842) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31960) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18999) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1982) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3174) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26043) * $signed(input_fmap_108[7:0]) +
	( 11'sd 972) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12984) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20113) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11023) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31743) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14986) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20696) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25262) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10173) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29124) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5835) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28675) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29319) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 16'sd 21106) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1627) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11712) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_6[7:0]) +
	( 9'sd 159) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32450) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28974) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16976) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3334) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5154) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18075) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26200) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31574) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20889) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9551) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23934) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29047) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7500) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14253) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24786) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3517) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9358) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25992) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17245) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16636) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14302) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_38[7:0]) +
	( 11'sd 766) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8497) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17053) * $signed(input_fmap_43[7:0]) +
	( 13'sd 4068) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18798) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14569) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23530) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5908) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25060) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17297) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13159) * $signed(input_fmap_55[7:0]) +
	( 10'sd 438) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5120) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21896) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21953) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30402) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14278) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8093) * $signed(input_fmap_65[7:0]) +
	( 11'sd 803) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9842) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10598) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25491) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18283) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6574) * $signed(input_fmap_74[7:0]) +
	( 12'sd 2039) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4878) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22752) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11312) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24341) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6026) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22200) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27265) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9341) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13753) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24369) * $signed(input_fmap_85[7:0]) +
	( 11'sd 796) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12736) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2322) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17680) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23901) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21703) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8107) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20529) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28857) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21189) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8427) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6640) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15759) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4229) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3248) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16211) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24137) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5357) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32333) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27326) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19979) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10502) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2868) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22171) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3708) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15117) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16684) * $signed(input_fmap_125[7:0]) +
	( 12'sd 2015) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5396) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 16'sd 20487) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3072) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32765) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32355) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10796) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21337) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31100) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16059) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17209) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5706) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20279) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13023) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18292) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7589) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6338) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11396) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28288) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8134) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2861) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18238) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15948) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31555) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27918) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28723) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18612) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15554) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10679) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29037) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3946) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10048) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5096) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30331) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7859) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1074) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5598) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9167) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7873) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11637) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1956) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4658) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15292) * $signed(input_fmap_58[7:0]) +
	( 11'sd 771) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30932) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26181) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30606) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16952) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16719) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16356) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13726) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21648) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23311) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27440) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24770) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32575) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13903) * $signed(input_fmap_84[7:0]) +
	( 10'sd 492) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17369) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10624) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5239) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32135) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24515) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24370) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3911) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29407) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29135) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28584) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21182) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18342) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23360) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26310) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13404) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18166) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20404) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5674) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29732) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8581) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3159) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25952) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13728) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26795) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13007) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25366) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 15'sd 10386) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32243) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19444) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_6[7:0]) +
	( 11'sd 777) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18058) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1446) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6918) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31445) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21796) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5562) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5627) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30739) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27454) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29941) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12733) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14553) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18173) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32379) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17115) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7515) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28272) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7434) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30560) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27526) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5198) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11224) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5124) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6847) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6761) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25881) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18188) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15388) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17458) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14520) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24642) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16926) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8066) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9155) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15261) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22003) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32235) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5595) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27710) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10508) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12810) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1727) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16333) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19907) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3229) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8970) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7835) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2250) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6617) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23240) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7565) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26846) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9987) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21489) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26268) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25298) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15103) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16077) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4149) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20076) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7379) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20034) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6627) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9030) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15751) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3709) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6264) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14008) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4591) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3206) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13743) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5248) * $signed(input_fmap_109[7:0]) +
	( 8'sd 107) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11442) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22324) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29891) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18725) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13627) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10056) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18085) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1654) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4981) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31681) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 15'sd 8839) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19459) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28714) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5918) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11981) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5668) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18114) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1132) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15844) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13075) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22707) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22543) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2524) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13892) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25205) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13486) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28204) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20334) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31620) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17326) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23988) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3442) * $signed(input_fmap_27[7:0]) +
	( 10'sd 371) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10517) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25448) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9436) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9502) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22372) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27860) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7166) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6458) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5197) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14591) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29338) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30859) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2506) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10307) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11722) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14990) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13708) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10857) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28285) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30466) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22950) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4780) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22323) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31701) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30468) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16682) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16659) * $signed(input_fmap_71[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11188) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22507) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32048) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9393) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12219) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17590) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29923) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4125) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25068) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3089) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4813) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17842) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21379) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19672) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29339) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3823) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15407) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6434) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12929) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29980) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14821) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14994) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8668) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28163) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20347) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11165) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32215) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20116) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4762) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6319) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5322) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18393) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15875) * $signed(input_fmap_124[7:0]) +
	( 11'sd 852) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29351) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 16'sd 24632) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13380) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9834) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20235) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28641) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24166) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2656) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22451) * $signed(input_fmap_10[7:0]) +
	( 11'sd 943) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27152) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10412) * $signed(input_fmap_14[7:0]) +
	( 11'sd 937) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17708) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13985) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4201) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5644) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7061) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7131) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16785) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11637) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28308) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10993) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11328) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27464) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4346) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31090) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30455) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12999) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27711) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4511) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28138) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26667) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26582) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30830) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18362) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15282) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2588) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11734) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17746) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18631) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23208) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31199) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21914) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16361) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_75[7:0]) +
	( 10'sd 357) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5302) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4384) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9144) * $signed(input_fmap_79[7:0]) +
	( 11'sd 578) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17331) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28705) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7446) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11396) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27641) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13852) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6385) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20087) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16712) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13051) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19069) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21725) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22342) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8972) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32043) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31192) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23147) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10074) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28747) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32493) * $signed(input_fmap_111[7:0]) +
	( 11'sd 695) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23616) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19519) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_116[7:0]) +
	( 10'sd 466) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8400) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3494) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31782) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30838) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9574) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15702) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9291) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 15'sd 9083) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19254) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11357) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30748) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2209) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4759) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8534) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13182) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_14[7:0]) +
	( 10'sd 322) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8093) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11286) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20482) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18772) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2854) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20846) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15328) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26429) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16145) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13194) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6204) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11597) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21277) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18955) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22710) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1762) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2697) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18167) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6627) * $signed(input_fmap_39[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14421) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15599) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10913) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2858) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16491) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32245) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18185) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6417) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31860) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10466) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23310) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19493) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26144) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1899) * $signed(input_fmap_71[7:0]) +
	( 14'sd 8091) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_73[7:0]) +
	( 11'sd 524) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31327) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20685) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24602) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32388) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22593) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21312) * $signed(input_fmap_85[7:0]) +
	( 11'sd 629) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15016) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27025) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17350) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6863) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16953) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30223) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26850) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14958) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24440) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29327) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5103) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21595) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6516) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13210) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9696) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18446) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28277) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10794) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1219) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9069) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10008) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23911) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8952) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7489) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9157) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19152) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11703) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 16'sd 19969) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6521) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11273) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9842) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19644) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17201) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4126) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12226) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27470) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15414) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29253) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14564) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16184) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_18[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2973) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9888) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17167) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18138) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12593) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20986) * $signed(input_fmap_26[7:0]) +
	( 10'sd 390) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8601) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11753) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21734) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5677) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4497) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1386) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22543) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8451) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6717) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11090) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29711) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14504) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32709) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15848) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17473) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17608) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8306) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12660) * $signed(input_fmap_63[7:0]) +
	( 11'sd 790) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2091) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14310) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9065) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18600) * $signed(input_fmap_68[7:0]) +
	( 9'sd 218) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27568) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29374) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5093) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28508) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13020) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28139) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5722) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26120) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5293) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23638) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15919) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24955) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26180) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24841) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25734) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21168) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2986) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22380) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29887) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9606) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29711) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31246) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14265) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19420) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14376) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20865) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8395) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14331) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7171) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6497) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8332) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8352) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1813) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31940) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13928) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9468) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2550) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10403) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31010) * $signed(input_fmap_124[7:0]) +
	( 11'sd 948) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25314) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 16'sd 24199) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17055) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8864) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4667) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15472) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16025) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16928) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10679) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10619) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10545) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12007) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8090) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25242) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3637) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20375) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5515) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10007) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26867) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23958) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31775) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15895) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8861) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14194) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17165) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17371) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11320) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24109) * $signed(input_fmap_34[7:0]) +
	( 10'sd 436) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1761) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1926) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10810) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25235) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_49[7:0]) +
	( 10'sd 361) * $signed(input_fmap_50[7:0]) +
	( 14'sd 8048) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7130) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2887) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32175) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29675) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6498) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17441) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6652) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15972) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13513) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19801) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3057) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12791) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2545) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18886) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5237) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29313) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6013) * $signed(input_fmap_78[7:0]) +
	( 9'sd 153) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25945) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14713) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6439) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18734) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8705) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6636) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2783) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20148) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10309) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12529) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20424) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2860) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9725) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17074) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14448) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20872) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26726) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23869) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1575) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21383) * $signed(input_fmap_108[7:0]) +
	( 7'sd 44) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10697) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13758) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15507) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7187) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32572) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24192) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29629) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7059) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32347) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31432) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6959) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 15'sd 15721) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31181) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16940) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21407) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22561) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18038) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10536) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_11[7:0]) +
	( 11'sd 600) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1828) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13416) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13433) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9403) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11580) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25819) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23771) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25621) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20918) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12992) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17583) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11995) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3597) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21520) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10698) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30181) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16793) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31164) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31349) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12566) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30043) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18638) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17159) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28264) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32400) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21648) * $signed(input_fmap_46[7:0]) +
	( 9'sd 206) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_48[7:0]) +
	( 13'sd 4004) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21811) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29996) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22465) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6013) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11646) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3115) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30659) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30406) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13504) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20295) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6698) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27651) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6678) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13792) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6491) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31833) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14369) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5162) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_77[7:0]) +
	( 11'sd 968) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9496) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2876) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30486) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10927) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26332) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5425) * $signed(input_fmap_88[7:0]) +
	( 10'sd 310) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18041) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28596) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27966) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22300) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24454) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5440) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24698) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27726) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5040) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4427) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11002) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23350) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27603) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28475) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27945) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7688) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22935) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13154) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4921) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1065) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7365) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28649) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17355) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13989) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3536) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27383) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 16'sd 22562) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3157) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1338) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18522) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18370) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7521) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27863) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1050) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15785) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12218) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8838) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3600) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7096) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27466) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32542) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29347) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2157) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27029) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5149) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20465) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17431) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27314) * $signed(input_fmap_35[7:0]) +
	( 11'sd 810) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2647) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21029) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27904) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17746) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12248) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6338) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23903) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18769) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3781) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1483) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7529) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31213) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16044) * $signed(input_fmap_54[7:0]) +
	( 11'sd 722) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8542) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31731) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21685) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28717) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31724) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2629) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9520) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24974) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27466) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4765) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6000) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27218) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22068) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13587) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13649) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11157) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30611) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28535) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18196) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7844) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1134) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20388) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21041) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27009) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7181) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19555) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26564) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2790) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12910) * $signed(input_fmap_95[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5159) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27332) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7609) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20936) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28331) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30949) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2955) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22892) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31419) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32441) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12243) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10299) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15168) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32601) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18577) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9099) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7799) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12177) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30646) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8635) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31881) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26731) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 16'sd 28515) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21045) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6381) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7051) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14569) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32426) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4751) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4343) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8228) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23116) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11550) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16043) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7204) * $signed(input_fmap_20[7:0]) +
	( 9'sd 172) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3077) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5024) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32639) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2694) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4909) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27479) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29799) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7352) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11346) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5950) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7018) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25086) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6374) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6207) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2123) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29868) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21818) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30380) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14185) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27833) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31635) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27468) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16897) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25669) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31499) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23180) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28287) * $signed(input_fmap_61[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25998) * $signed(input_fmap_63[7:0]) +
	( 11'sd 788) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2595) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30368) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24373) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23251) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18430) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18770) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22512) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15092) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10078) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16828) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14182) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10803) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20940) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20317) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18838) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9712) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_88[7:0]) +
	( 7'sd 46) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24513) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9302) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27543) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28651) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11570) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12326) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32296) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16225) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25370) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14250) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24157) * $signed(input_fmap_104[7:0]) +
	( 7'sd 42) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22058) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25111) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31041) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_110[7:0]) +
	( 9'sd 162) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11214) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25230) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3950) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_119[7:0]) +
	( 11'sd 591) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9351) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21967) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3349) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13634) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6675) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 16'sd 17086) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12812) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6524) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24188) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1221) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20798) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2490) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4957) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21177) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26714) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22382) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26973) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9234) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26420) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8982) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10979) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20950) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9395) * $signed(input_fmap_26[7:0]) +
	( 10'sd 385) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28553) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12970) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26736) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32533) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2506) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10327) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8815) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32743) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2933) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31426) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11095) * $signed(input_fmap_46[7:0]) +
	( 10'sd 301) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9304) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14450) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30609) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28098) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27093) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30189) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22523) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5962) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22471) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21949) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28405) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12991) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11822) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19885) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11808) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21679) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8986) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28888) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25233) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29994) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5069) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24436) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26944) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7968) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12191) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20717) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31249) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11945) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28692) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23457) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12931) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29686) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28102) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16800) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27518) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22784) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24280) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14837) * $signed(input_fmap_105[7:0]) +
	( 10'sd 472) * $signed(input_fmap_106[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21856) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6334) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3768) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5573) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29043) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30575) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15632) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28697) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3676) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1337) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25936) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 16'sd 28566) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8218) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20632) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12704) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24422) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31063) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19244) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31288) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25177) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32443) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30251) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8112) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7201) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4188) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15283) * $signed(input_fmap_19[7:0]) +
	( 11'sd 590) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25230) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_22[7:0]) +
	( 13'sd 4018) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22000) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20195) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19290) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15111) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6511) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22764) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14872) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26141) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7130) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22163) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6520) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14347) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19667) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15191) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21007) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2483) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11192) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13055) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32273) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28411) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12083) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22297) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21829) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3566) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16083) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5426) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14901) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14045) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23973) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6498) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16270) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13618) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12268) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22558) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20691) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10263) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18650) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6663) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12161) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1422) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13020) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30553) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11107) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13065) * $signed(input_fmap_86[7:0]) +
	( 14'sd 8067) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7679) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25780) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24121) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25131) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7637) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4653) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20969) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30779) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23755) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7277) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15164) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20669) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16473) * $signed(input_fmap_110[7:0]) +
	( 15'sd 16247) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32662) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14384) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10086) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1755) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29613) * $signed(input_fmap_123[7:0]) +
	( 9'sd 173) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3600) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8344) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32466) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 16'sd 29666) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6658) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4933) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11960) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5710) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22854) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8265) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1164) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7926) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3935) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26660) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14195) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24751) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5336) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18683) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18873) * $signed(input_fmap_24[7:0]) +
	( 10'sd 373) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27799) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32590) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3035) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13672) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27406) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7552) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23946) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17546) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30910) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2089) * $signed(input_fmap_43[7:0]) +
	( 9'sd 150) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3195) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23072) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15140) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3880) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11250) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30089) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1791) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17612) * $signed(input_fmap_57[7:0]) +
	( 10'sd 265) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27710) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13123) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14873) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18589) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28160) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2671) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7968) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12636) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9752) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13404) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24703) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20564) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29805) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28470) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19947) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28033) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4676) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3783) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30106) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22932) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28288) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21174) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7308) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6536) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28058) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9921) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26817) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29556) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18702) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13113) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15263) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11859) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21354) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19746) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7215) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_113[7:0]) +
	( 7'sd 48) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15713) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2233) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_121[7:0]) +
	( 10'sd 294) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19996) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11207) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11515) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19706) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 16'sd 17080) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24285) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10271) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16991) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12021) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10645) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19534) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2943) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16720) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26664) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22632) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11666) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22564) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17211) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16192) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17355) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26789) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31152) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20233) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14956) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17798) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3274) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9804) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8200) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7767) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15112) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12791) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12428) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19468) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9889) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2794) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18062) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28548) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27064) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17542) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28294) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2836) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22069) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8760) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20206) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5052) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14408) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26340) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25998) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1158) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25748) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19935) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4243) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32675) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9055) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21613) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17677) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2318) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11189) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20352) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27733) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24137) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26524) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27499) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19897) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11814) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5990) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32574) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6811) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14669) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23710) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2113) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8780) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23574) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31741) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31590) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2229) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27607) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17026) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30431) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9856) * $signed(input_fmap_99[7:0]) +
	( 11'sd 768) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12410) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32663) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3305) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15624) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8171) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7615) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31713) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21884) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5120) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30816) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32357) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16235) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27409) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26382) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14133) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3512) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 16'sd 22750) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30896) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4883) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19458) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6925) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19556) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2505) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30197) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18053) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32235) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1381) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13800) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8595) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10692) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5932) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17851) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16024) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24308) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11702) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15847) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16725) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15971) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24614) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21675) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30382) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15987) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16821) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5216) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14398) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8323) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29698) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11778) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1332) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1291) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24644) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3488) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21709) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6338) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25531) * $signed(input_fmap_67[7:0]) +
	( 14'sd 8096) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4775) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24063) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20711) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16807) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31271) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16234) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10745) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11784) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30321) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4428) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29303) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_82[7:0]) +
	( 9'sd 248) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_84[7:0]) +
	( 11'sd 516) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14105) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4272) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15101) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8459) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3205) * $signed(input_fmap_93[7:0]) +
	( 11'sd 877) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30715) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18767) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16949) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19830) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31600) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20659) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9002) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18867) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27456) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15282) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31313) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8882) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1449) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_112[7:0]) +
	( 10'sd 464) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1546) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5263) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30162) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31679) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7579) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11988) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6934) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5827) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2067) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 14'sd 8067) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17959) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6790) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26152) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3442) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5847) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14665) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18535) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3120) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20573) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5055) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21905) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6931) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17186) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28220) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9246) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18053) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17267) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6136) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14764) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7278) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17511) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20441) * $signed(input_fmap_29[7:0]) +
	( 14'sd 8032) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30253) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22936) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14074) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6039) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29983) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26098) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12462) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27729) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28367) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32366) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23473) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26737) * $signed(input_fmap_48[7:0]) +
	( 6'sd 26) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23798) * $signed(input_fmap_51[7:0]) +
	( 11'sd 757) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9565) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30532) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19385) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6862) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3365) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20996) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6552) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5459) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18954) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19251) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26053) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20356) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25475) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22175) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25512) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_72[7:0]) +
	( 10'sd 264) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18487) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25662) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16483) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26200) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18989) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31891) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22114) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19556) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16020) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16049) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27428) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4765) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28128) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4236) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21406) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26788) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3926) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11785) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5714) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11934) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20655) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30015) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4507) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9297) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4332) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12255) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29291) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19349) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17100) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17826) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7104) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14010) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12508) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31867) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31648) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32197) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6206) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15216) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1935) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2081) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 15'sd 8370) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3990) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17928) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3110) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19876) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9861) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26532) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_11[7:0]) +
	( 11'sd 989) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25085) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10381) * $signed(input_fmap_14[7:0]) +
	( 14'sd 8153) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4571) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21437) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15393) * $signed(input_fmap_22[7:0]) +
	( 10'sd 330) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28535) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21283) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31380) * $signed(input_fmap_27[7:0]) +
	( 11'sd 968) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30712) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27645) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12226) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15754) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32162) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10461) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6576) * $signed(input_fmap_38[7:0]) +
	( 14'sd 8067) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29332) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11133) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2452) * $signed(input_fmap_49[7:0]) +
	( 10'sd 363) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23116) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16514) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32048) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_56[7:0]) +
	( 11'sd 533) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13105) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2961) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29858) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18125) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8763) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24007) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6024) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32091) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7469) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1746) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9461) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7098) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18858) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15364) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4499) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14886) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20372) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1073) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14097) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28563) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6362) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9526) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28831) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6095) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6274) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10471) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19925) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6540) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23701) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16933) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14828) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3003) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19653) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7712) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9232) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14236) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15515) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1447) * $signed(input_fmap_117[7:0]) +
	( 13'sd 4040) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11210) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24018) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2131) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14346) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12481) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12525) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 16'sd 24202) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13561) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5111) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20102) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24071) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6158) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24158) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16373) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25022) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21177) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11287) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22015) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1433) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5576) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12890) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13182) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10715) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26708) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29081) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4875) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22703) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28866) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1727) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16669) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21090) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17267) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31277) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8593) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5641) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19269) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18990) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14491) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6502) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_58[7:0]) +
	( 12'sd 2001) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32191) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15807) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16336) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6788) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25435) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4622) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30457) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30919) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17375) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31650) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32747) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24569) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5968) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12648) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27549) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28517) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14837) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20450) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15289) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9516) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29474) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12428) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14269) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9808) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4374) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_103[7:0]) +
	( 11'sd 745) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12968) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24781) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27556) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23210) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24328) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1885) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12123) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3426) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19036) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29947) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9606) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9791) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12320) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9071) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6522) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 14'sd 5719) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12161) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20741) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30437) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24542) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3721) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13307) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16867) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17488) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_11[7:0]) +
	( 11'sd 736) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23517) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19625) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16247) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2243) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22268) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18564) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13164) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10702) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4700) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1700) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10134) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2768) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9121) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12866) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9965) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25859) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1605) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14471) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30319) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8664) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20507) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12766) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2299) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10539) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1832) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23969) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29101) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11641) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7923) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6561) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6420) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10533) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29492) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8362) * $signed(input_fmap_70[7:0]) +
	( 11'sd 975) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26962) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7935) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5736) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15783) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2124) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29402) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7837) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30193) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27437) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31847) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12867) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28787) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_88[7:0]) +
	( 11'sd 662) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2377) * $signed(input_fmap_90[7:0]) +
	( 14'sd 8000) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27418) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31357) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24549) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9229) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28006) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12212) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18052) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25906) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24633) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6948) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25969) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31334) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15472) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27347) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25516) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16998) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10269) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20055) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15591) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26906) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 16'sd 23102) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6595) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32005) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2927) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20687) * $signed(input_fmap_4[7:0]) +
	( 11'sd 980) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7249) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30698) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14797) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9758) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12249) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27132) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17802) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6331) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27533) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23687) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5348) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1422) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31280) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18609) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7483) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23371) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9679) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9575) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2367) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13495) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21941) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11047) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21052) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20571) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19584) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11724) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_43[7:0]) +
	( 3'sd 3) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25396) * $signed(input_fmap_45[7:0]) +
	( 11'sd 696) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23697) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18276) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15981) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23356) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_56[7:0]) +
	( 11'sd 847) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19103) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25751) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30362) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17085) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24479) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24341) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32593) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14027) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10827) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30948) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6222) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5574) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20001) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27662) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6788) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25652) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4179) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26781) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31733) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10405) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21072) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27921) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28730) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20096) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22343) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14896) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9436) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19603) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2159) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5887) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23039) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30944) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1512) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31285) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20135) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_107[7:0]) +
	( 11'sd 1019) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8362) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9852) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18913) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4193) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12953) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24562) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24578) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 16'sd 24097) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26885) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29140) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4992) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20566) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1083) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3358) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26572) * $signed(input_fmap_15[7:0]) +
	( 7'sd 61) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20227) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24819) * $signed(input_fmap_20[7:0]) +
	( 9'sd 153) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9099) * $signed(input_fmap_22[7:0]) +
	( 11'sd 533) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21877) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8809) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20660) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31238) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29753) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14371) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15725) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30289) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31722) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30264) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23675) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13078) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31534) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6503) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16197) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2553) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4958) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7460) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32751) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9944) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6168) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1041) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6068) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2512) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22665) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5381) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14671) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31705) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24739) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30189) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14057) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24312) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11001) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30277) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14156) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6631) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13426) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32580) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3421) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26469) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12856) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7943) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10244) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25116) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11734) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_114[7:0]) +
	( 10'sd 383) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13872) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23252) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26707) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23166) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28025) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27636) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31621) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25258) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 15'sd 12824) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1817) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29072) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6375) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25323) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19421) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14460) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19834) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1363) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31497) * $signed(input_fmap_11[7:0]) +
	( 11'sd 618) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25503) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14008) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10612) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27471) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16969) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8749) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16170) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9885) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25260) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18420) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19591) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21616) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5328) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31808) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12884) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4690) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23335) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14863) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12836) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17018) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9705) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5211) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31857) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15248) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2502) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31684) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30127) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14610) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27264) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2236) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32153) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32510) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9265) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28466) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2239) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28980) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8512) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14874) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8603) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31244) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14864) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5423) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24094) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26054) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27284) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7522) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9244) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12299) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30714) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31498) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28668) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23412) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3285) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32453) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10607) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4978) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32291) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18540) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13344) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8011) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10552) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14089) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21359) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20767) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4776) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23503) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2533) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10283) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9952) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26254) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11664) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27427) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18223) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 26783) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6864) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10075) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17945) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21831) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24071) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29859) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29503) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25778) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12214) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8148) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6751) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21960) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27365) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21491) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5593) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7884) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7029) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11890) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19506) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10271) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5418) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12233) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14781) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16401) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22102) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2631) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1865) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24886) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3694) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19647) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13553) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18168) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18123) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12366) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26943) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4773) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15877) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22129) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_61[7:0]) +
	( 13'sd 4042) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7667) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27985) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9937) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7166) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1118) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23299) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19345) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10490) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3726) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1193) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14604) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17490) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20857) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25123) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7831) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27442) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25813) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_93[7:0]) +
	( 10'sd 312) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20570) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1116) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17600) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23257) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26858) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1846) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17758) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3142) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7118) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15158) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15246) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30504) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2856) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16339) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32691) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31444) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18904) * $signed(input_fmap_121[7:0]) +
	( 10'sd 373) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19521) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10061) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16183) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 16'sd 29448) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25305) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31698) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26849) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27292) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1737) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30869) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8063) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23533) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15638) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21412) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7804) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24611) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32684) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28594) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32383) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5618) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17021) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30831) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9194) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3099) * $signed(input_fmap_24[7:0]) +
	( 11'sd 707) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15447) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15595) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26503) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29633) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_34[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22448) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2493) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28141) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16812) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30497) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5796) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7826) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16544) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1912) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16645) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15538) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2967) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26762) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5527) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24860) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9896) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31909) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19578) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22744) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8295) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15772) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29765) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30242) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24358) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9414) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24750) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9536) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3269) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28780) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24337) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28538) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11584) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4728) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12609) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8825) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23053) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29082) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18554) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12284) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27321) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10086) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19155) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3601) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8980) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1547) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27528) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4735) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2498) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13937) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6356) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13285) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19830) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24742) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20939) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11291) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29608) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26509) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_123[7:0]) +
	( 11'sd 558) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10221) * $signed(input_fmap_125[7:0]) +
	( 9'sd 184) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16314) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 14'sd 5949) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32068) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20294) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3824) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4871) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27997) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13229) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25909) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17949) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1612) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21788) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31353) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24578) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26063) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2795) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2710) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23555) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31351) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14478) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2730) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26001) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10526) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32494) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17957) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10362) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13128) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21638) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15190) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5375) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24239) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5429) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_55[7:0]) +
	( 7'sd 56) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31506) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8635) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22325) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15518) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30758) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7966) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2644) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2107) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6306) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9891) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9691) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11441) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28046) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24222) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16872) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5738) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26382) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14771) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5822) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25982) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32692) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2432) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28866) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12268) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10722) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16466) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31620) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10118) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15293) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13887) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20617) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10757) * $signed(input_fmap_108[7:0]) +
	( 11'sd 890) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9063) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13134) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14473) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4384) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28427) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1740) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14502) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5710) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13421) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19869) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25465) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 16'sd 32306) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5340) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1714) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18119) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30709) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23883) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7963) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29898) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30789) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7240) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15355) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7114) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20253) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14631) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21896) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21220) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21160) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25478) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24826) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3141) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11703) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31463) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15695) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15387) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20289) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9183) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24913) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20908) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5898) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10009) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15789) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25478) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27660) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14955) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31062) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23905) * $signed(input_fmap_61[7:0]) +
	( 11'sd 620) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14582) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30617) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9337) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24613) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23841) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24169) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17642) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18256) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7320) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21327) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19502) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5718) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13938) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7963) * $signed(input_fmap_81[7:0]) +
	( 10'sd 330) * $signed(input_fmap_82[7:0]) +
	( 11'sd 874) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27034) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5914) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25805) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8856) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16629) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21562) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18597) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17216) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2766) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3410) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21580) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4578) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6722) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26321) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32682) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30036) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12049) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1635) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1028) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3728) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23844) * $signed(input_fmap_112[7:0]) +
	( 12'sd 2025) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11003) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16078) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6060) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4418) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7092) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25239) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9932) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18361) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27066) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3872) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9776) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 15'sd 13249) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17873) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5988) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32535) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8209) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8042) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14870) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7749) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26040) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9342) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12219) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3340) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26844) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14718) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23486) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2652) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2588) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5378) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28643) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6049) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21688) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3133) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14644) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26574) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21003) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8262) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20770) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14286) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1350) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21347) * $signed(input_fmap_41[7:0]) +
	( 9'sd 255) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27580) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8260) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28933) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10721) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26360) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31448) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19110) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6194) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24566) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7650) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7358) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3114) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25168) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1231) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26088) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20758) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1383) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18043) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24422) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29906) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22478) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_73[7:0]) +
	( 14'sd 8155) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12087) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18051) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25781) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31670) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26314) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2485) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31732) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2427) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21704) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27210) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22133) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24648) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3094) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13594) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21008) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3236) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30575) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10993) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4653) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29482) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26801) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3620) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8564) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31391) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27064) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17493) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16503) * $signed(input_fmap_124[7:0]) +
	( 11'sd 977) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5531) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28712) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 16'sd 26714) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22495) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15206) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14348) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9327) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12798) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9940) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4404) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31746) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21939) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6969) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8466) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26183) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15776) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32553) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31419) * $signed(input_fmap_20[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5458) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32187) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6105) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25916) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17128) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12079) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8315) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28215) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25143) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13349) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10340) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29101) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21388) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25253) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10841) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19060) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12764) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17788) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4376) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21626) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8649) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1179) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1915) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25239) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11471) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25153) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_60[7:0]) +
	( 11'sd 571) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24801) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15137) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30844) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3559) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11758) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14297) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13619) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30058) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24142) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32577) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21894) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17181) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27634) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24638) * $signed(input_fmap_81[7:0]) +
	( 8'sd 78) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27374) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19054) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30397) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16233) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8431) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13029) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27206) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18262) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22407) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30529) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26656) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32214) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23731) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8554) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23582) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17333) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12505) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5217) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_110[7:0]) +
	( 9'sd 131) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6215) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31653) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_116[7:0]) +
	( 10'sd 370) * $signed(input_fmap_117[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13695) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_122[7:0]) +
	( 11'sd 589) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9527) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 16'sd 27429) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22702) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11407) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25294) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15688) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12465) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10049) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31944) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25662) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28706) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31056) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22761) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14099) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12135) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1712) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9450) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24180) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6134) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21014) * $signed(input_fmap_26[7:0]) +
	( 9'sd 176) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26448) * $signed(input_fmap_30[7:0]) +
	( 11'sd 839) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11310) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29540) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31919) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12452) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8820) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12433) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27112) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7737) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19007) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23963) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22255) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9008) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13886) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24408) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_54[7:0]) +
	( 13'sd 4004) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21717) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22964) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2118) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18543) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27749) * $signed(input_fmap_60[7:0]) +
	( 11'sd 996) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12547) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6905) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9492) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24970) * $signed(input_fmap_66[7:0]) +
	( 6'sd 26) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3157) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13439) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21201) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21661) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1347) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_76[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30961) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_79[7:0]) +
	( 11'sd 786) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30954) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11011) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20059) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2556) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26895) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16922) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18688) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31361) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28875) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22237) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13749) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26132) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27490) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30489) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25250) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29834) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5474) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1098) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6923) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10319) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20661) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32051) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15358) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_112[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7755) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24921) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31782) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15539) * $signed(input_fmap_119[7:0]) +
	( 11'sd 581) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16293) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30613) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26579) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21729) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18120) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8872) * $signed(input_fmap_126[7:0]) +
	( 11'sd 907) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 16'sd 25293) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1554) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9141) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26566) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5090) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30154) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14682) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16432) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16215) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16062) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24697) * $signed(input_fmap_11[7:0]) +
	( 9'sd 152) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22203) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22380) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8016) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20565) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16361) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19609) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1314) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23552) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8601) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24560) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9311) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16081) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15795) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30115) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8418) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2250) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30501) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27665) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15814) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11411) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11390) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19589) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14230) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9371) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28150) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20741) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10650) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3948) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8637) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5457) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6365) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3788) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24503) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8537) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6946) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22645) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13734) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1915) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3822) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31247) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3478) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25022) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26935) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26664) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23042) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29469) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31146) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32724) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15042) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10800) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29278) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3400) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24425) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24782) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19406) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23792) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29231) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9568) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19057) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23766) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3413) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25564) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11061) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32584) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13475) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17608) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21279) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23326) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17640) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4980) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30045) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30154) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 16'sd 21918) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30691) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_6[7:0]) +
	( 10'sd 412) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18729) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3969) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8787) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_13[7:0]) +
	( 14'sd 8097) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23124) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28956) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29786) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8651) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30345) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24909) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26512) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11595) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14576) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20244) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13468) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4692) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21148) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9803) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4643) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19679) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3873) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12090) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2186) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1994) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2746) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17996) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6458) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10726) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32226) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25788) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4373) * $signed(input_fmap_61[7:0]) +
	( 11'sd 775) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15886) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15956) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4749) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11086) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32057) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30136) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21032) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31798) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10409) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23279) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28884) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20668) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_77[7:0]) +
	( 14'sd 8128) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19218) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21713) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1661) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10514) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11324) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29188) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31639) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24786) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31399) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14008) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15040) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31177) * $signed(input_fmap_94[7:0]) +
	( 11'sd 799) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14664) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12694) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22055) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5021) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11013) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7457) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32102) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10171) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27710) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7432) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25094) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27467) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28060) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10431) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21291) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4584) * $signed(input_fmap_117[7:0]) +
	( 10'sd 443) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29884) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_120[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16734) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16258) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18774) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 14'sd 6159) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26304) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21464) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2657) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1285) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21431) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3584) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21335) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_14[7:0]) +
	( 13'sd 4009) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21169) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4288) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10646) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18328) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22632) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28433) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13146) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6503) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3944) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32147) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30098) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14659) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5175) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19723) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21664) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3155) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23517) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30601) * $signed(input_fmap_36[7:0]) +
	( 11'sd 972) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29537) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8812) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21888) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5093) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8138) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32512) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21910) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17815) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7398) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27001) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1644) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16236) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4655) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13098) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2701) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15670) * $signed(input_fmap_72[7:0]) +
	( 6'sd 27) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14287) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10431) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30957) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9315) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16602) * $signed(input_fmap_80[7:0]) +
	( 9'sd 159) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31826) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6316) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24151) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26839) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26927) * $signed(input_fmap_89[7:0]) +
	( 10'sd 353) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25875) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32143) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17499) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23095) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16834) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29343) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6510) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15225) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23662) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28833) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23784) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27385) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6346) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6933) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16968) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1649) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15604) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23607) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30769) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2722) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_123[7:0]) +
	( 11'sd 874) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17227) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22087) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 13'sd 2658) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17863) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25435) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11465) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27135) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9836) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12663) * $signed(input_fmap_12[7:0]) +
	( 14'sd 8173) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3773) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3407) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21726) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22288) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19016) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1524) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20652) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10450) * $signed(input_fmap_22[7:0]) +
	( 11'sd 758) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5709) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23993) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13505) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27218) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4479) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4122) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23486) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2709) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29016) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25446) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14546) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25536) * $signed(input_fmap_44[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18736) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8780) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27232) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30381) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2250) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28716) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7181) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12087) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18719) * $signed(input_fmap_58[7:0]) +
	( 12'sd 2000) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13480) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13594) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22168) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27822) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9821) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2451) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18890) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15978) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21967) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23265) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1318) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2827) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3386) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2743) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7886) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4100) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29001) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2729) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7370) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27765) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8555) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29438) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9965) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_110[7:0]) +
	( 9'sd 149) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18837) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28983) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2835) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_122[7:0]) +
	( 8'sd 74) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_124[7:0]) +
	( 11'sd 991) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4311) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 16'sd 23087) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32586) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17500) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32705) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24542) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15680) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14287) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2182) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11612) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10804) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30781) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20642) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13918) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7523) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19769) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11997) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5028) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16666) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13465) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7199) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24024) * $signed(input_fmap_30[7:0]) +
	( 11'sd 875) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1418) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25278) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5055) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14588) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20720) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26224) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_40[7:0]) +
	( 11'sd 673) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25272) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2493) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22728) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5716) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5815) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29538) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25774) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17641) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10813) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16097) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6591) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13905) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28643) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_60[7:0]) +
	( 10'sd 354) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18165) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30704) * $signed(input_fmap_63[7:0]) +
	( 11'sd 930) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16856) * $signed(input_fmap_65[7:0]) +
	( 11'sd 847) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27732) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6827) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2124) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19039) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9746) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3328) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29987) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14650) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17090) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28528) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14082) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27427) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7276) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3543) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11444) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32709) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6653) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32273) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30546) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29972) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10583) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24701) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31926) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19850) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6822) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32353) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30059) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1712) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13497) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25320) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15533) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18947) * $signed(input_fmap_123[7:0]) +
	( 10'sd 288) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11253) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31480) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 16'sd 24759) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28798) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29261) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1664) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14435) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27828) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17001) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_9[7:0]) +
	( 8'sd 83) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15008) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18109) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20211) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28739) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7491) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17378) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15916) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12016) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30961) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3494) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_36[7:0]) +
	( 10'sd 382) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8590) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21604) * $signed(input_fmap_39[7:0]) +
	( 8'sd 107) * $signed(input_fmap_40[7:0]) +
	( 11'sd 865) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6895) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23168) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27868) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17521) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25759) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18649) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16439) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27948) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31769) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15314) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5432) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7005) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_60[7:0]) +
	( 11'sd 780) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13071) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8333) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3414) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18074) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26449) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11982) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19544) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18835) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10770) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17260) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11933) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20084) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30813) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28773) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7583) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14134) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17354) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15430) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4937) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4117) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24870) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12573) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9387) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7612) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2655) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31918) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9731) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5176) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6568) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25080) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30737) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26074) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8059) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31397) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9244) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14254) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7693) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31869) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25562) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8867) * $signed(input_fmap_121[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21537) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10217) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 16'sd 26009) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4123) * $signed(input_fmap_1[7:0]) +
	( 11'sd 628) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3887) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1958) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28939) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8587) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25714) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3510) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14470) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7223) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10714) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20761) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14147) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3411) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19636) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_29[7:0]) +
	( 10'sd 486) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8892) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9034) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23584) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22929) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3581) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19180) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29053) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11007) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8242) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21463) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7828) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3585) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9246) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9618) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30753) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12124) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15134) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14819) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7530) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8628) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3761) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31733) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_63[7:0]) +
	( 7'sd 48) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31096) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7074) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30950) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23238) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5152) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13869) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7937) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6140) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10330) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23901) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31106) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21362) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9662) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21929) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31963) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26149) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13013) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10734) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15582) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2229) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13394) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19798) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1343) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15970) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2701) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3366) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10947) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17160) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2379) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14164) * $signed(input_fmap_118[7:0]) +
	( 10'sd 365) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6773) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25987) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19740) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4970) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20466) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32750) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 15'sd 15816) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25116) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11187) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18132) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3936) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2452) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17838) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1996) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22433) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27867) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9491) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2601) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22338) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23506) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27102) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32510) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16934) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25321) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24942) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8828) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3666) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32305) * $signed(input_fmap_34[7:0]) +
	( 11'sd 729) * $signed(input_fmap_35[7:0]) +
	( 7'sd 54) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12049) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3085) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5704) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5284) * $signed(input_fmap_41[7:0]) +
	( 9'sd 160) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29252) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1261) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9501) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32537) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19609) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27184) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9966) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20597) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8907) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9841) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24920) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21539) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10128) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1790) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3401) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27649) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29740) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29608) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15040) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5118) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12947) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29056) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22359) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20261) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17775) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24309) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9082) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14716) * $signed(input_fmap_84[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25874) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24465) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23544) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32197) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14798) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27444) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10252) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20485) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_96[7:0]) +
	( 11'sd 708) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22775) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6232) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20178) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27783) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25496) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2253) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5184) * $signed(input_fmap_108[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26250) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23760) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7328) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6891) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9473) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9384) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29599) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28610) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23833) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26060) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 16'sd 17282) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16411) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17227) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25738) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25040) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24050) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9781) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19900) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23148) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1536) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23214) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10669) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19698) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32510) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9877) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15796) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5399) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15440) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20348) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20377) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19558) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6590) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31764) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16110) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25160) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30428) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26424) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19294) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28917) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26737) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16055) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30033) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28298) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24928) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32519) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1332) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31076) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12199) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13152) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3493) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14299) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29299) * $signed(input_fmap_66[7:0]) +
	( 11'sd 739) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8470) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31814) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26758) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30056) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17867) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5768) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5964) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16839) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28905) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30876) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23167) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5303) * $signed(input_fmap_83[7:0]) +
	( 9'sd 212) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21489) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13644) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21652) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23787) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31670) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12643) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13660) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31630) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10070) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22733) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6497) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26741) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30382) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31897) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8831) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8598) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15522) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9182) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23026) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30298) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19370) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17730) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31493) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17379) * $signed(input_fmap_121[7:0]) +
	( 11'sd 1020) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2855) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17194) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 15'sd 11374) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4670) * $signed(input_fmap_1[7:0]) +
	( 11'sd 753) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6307) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5538) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14297) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15538) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21962) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23118) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28016) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26714) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29184) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21702) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5717) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1992) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19443) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10459) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4361) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10749) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7278) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26441) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23258) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5607) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24009) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28800) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6478) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24034) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9336) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14234) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1270) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11973) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23954) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13970) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12148) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26258) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9511) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32594) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10252) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24683) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24982) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22913) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17438) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9175) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21681) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14510) * $signed(input_fmap_69[7:0]) +
	( 11'sd 572) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15297) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1546) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23662) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18236) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31083) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3721) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7965) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15105) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31917) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10482) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19406) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24615) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17151) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19511) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3359) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19686) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7200) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21087) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23322) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17491) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15268) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5910) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4345) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9499) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31862) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16034) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6330) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13800) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13963) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8555) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5400) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15872) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22195) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1302) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12612) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8637) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10284) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23890) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9136) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26549) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2982) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23851) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14893) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17347) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 13'sd 2914) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24445) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22183) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19427) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4850) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18504) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26837) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_20[7:0]) +
	( 11'sd 1021) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12149) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20671) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13469) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18268) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6126) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13389) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16337) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28148) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7389) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26233) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32255) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10721) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18885) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18694) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9103) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7946) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19487) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24995) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23431) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19127) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9359) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2376) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5321) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15341) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30520) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10053) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21612) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15627) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22584) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19879) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20101) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21838) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9168) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5308) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24343) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26700) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11123) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6852) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19730) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24450) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3911) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18170) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14839) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11403) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25507) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21588) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11888) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31357) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9321) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30915) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15677) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18725) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24101) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22248) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8772) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19918) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28780) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4687) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3524) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28507) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6362) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25983) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22014) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 16'sd 27238) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12446) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20221) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9498) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22059) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5860) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11310) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20025) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2591) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19296) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32665) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11233) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6235) * $signed(input_fmap_20[7:0]) +
	( 9'sd 130) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17136) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25497) * $signed(input_fmap_25[7:0]) +
	( 11'sd 667) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16684) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29408) * $signed(input_fmap_29[7:0]) +
	( 6'sd 25) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20178) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28334) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28390) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10656) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30310) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4595) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11650) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4899) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21772) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7951) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10017) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26629) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21822) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15822) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17996) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12059) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21463) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29424) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20350) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31667) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6597) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13920) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6279) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24612) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25673) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11265) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8868) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27736) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32350) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22806) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24436) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2663) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31222) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2503) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30995) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23410) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20952) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5965) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10149) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28416) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8635) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14465) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9902) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3282) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21951) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2121) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8273) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15481) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8653) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11325) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13405) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14057) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22155) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17595) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27487) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31335) * $signed(input_fmap_121[7:0]) +
	( 10'sd 401) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1719) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28770) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28753) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11640) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 16'sd 25435) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24569) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32194) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14597) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21638) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_10[7:0]) +
	( 10'sd 475) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25399) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29067) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19420) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17332) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20821) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21661) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32449) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7165) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18378) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2556) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1874) * $signed(input_fmap_31[7:0]) +
	( 11'sd 937) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27373) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13870) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11904) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15514) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26893) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31769) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12672) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3225) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19136) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23410) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6837) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28954) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26397) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8073) * $signed(input_fmap_57[7:0]) +
	( 13'sd 4010) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24824) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32736) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24337) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16992) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23049) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28616) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26032) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_74[7:0]) +
	( 11'sd 594) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24159) * $signed(input_fmap_76[7:0]) +
	( 11'sd 955) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23509) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1238) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12244) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1408) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16916) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17453) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9343) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9408) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1865) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22916) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4922) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14481) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16611) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30368) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32420) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11802) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7403) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29966) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9911) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14225) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_102[7:0]) +
	( 9'sd 197) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10848) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25049) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26281) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1620) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12899) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8438) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5961) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29080) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11925) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32689) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 16'sd 31917) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10740) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15576) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10364) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7211) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17273) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8030) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23642) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10035) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16808) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18486) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21434) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1318) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24908) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11180) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4397) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19647) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32152) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17781) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5119) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20060) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10552) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15931) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13558) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3073) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12859) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8383) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30291) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25133) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16223) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10796) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21204) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15697) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22249) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28909) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16163) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5051) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26954) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11842) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14404) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17179) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21217) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16371) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31577) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8379) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5208) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17651) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28556) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1539) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21341) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3906) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3843) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12313) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28755) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19138) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19162) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14877) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30652) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21270) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23408) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31681) * $signed(input_fmap_83[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11065) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8285) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24147) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9024) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14693) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14057) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9647) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11760) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21664) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4893) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14789) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17095) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9876) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21004) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13590) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23875) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4192) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21014) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21326) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2920) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14117) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17307) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9464) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2984) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11426) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23117) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13217) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27562) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19685) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30114) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 15'sd 15748) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14274) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19162) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19742) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22717) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27244) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11924) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30506) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6205) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32651) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30820) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4453) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12110) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11054) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32748) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14284) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23569) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7476) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19295) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32553) * $signed(input_fmap_29[7:0]) +
	( 7'sd 62) * $signed(input_fmap_30[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2293) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31619) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20598) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23157) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14122) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29592) * $signed(input_fmap_40[7:0]) +
	( 11'sd 566) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8642) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6414) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23190) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6303) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26785) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20779) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4124) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29316) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12300) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25409) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27621) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29810) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15839) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19529) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3601) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11860) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19642) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12908) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30149) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1144) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3871) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12659) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9291) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31426) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19289) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28372) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16089) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18290) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32431) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26708) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32426) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30368) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5961) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17493) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22853) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15770) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24775) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8660) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1598) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26004) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16375) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29166) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22061) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19999) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32332) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_113[7:0]) +
	( 7'sd 55) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6869) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10325) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7213) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30339) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1535) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14200) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14306) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 15'sd 11819) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23669) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17862) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7818) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15321) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11632) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7535) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17791) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8236) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11712) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26753) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9226) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3042) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24031) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24868) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12682) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15016) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16283) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_27[7:0]) +
	( 10'sd 443) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6313) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1899) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3166) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16763) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2456) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3171) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26529) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11946) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16925) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26950) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_44[7:0]) +
	( 11'sd 675) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15605) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1101) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20037) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28458) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16543) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1536) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19570) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28420) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3606) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22175) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18340) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18862) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11337) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19914) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1992) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26126) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4993) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27873) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21885) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16307) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13378) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4328) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4446) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20111) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16142) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17312) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9395) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4236) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15598) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31409) * $signed(input_fmap_101[7:0]) +
	( 11'sd 780) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17639) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30886) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30786) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22252) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18688) * $signed(input_fmap_111[7:0]) +
	( 11'sd 851) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8878) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13544) * $signed(input_fmap_116[7:0]) +
	( 10'sd 409) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24813) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14672) * $signed(input_fmap_119[7:0]) +
	( 6'sd 30) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21513) * $signed(input_fmap_121[7:0]) +
	( 9'sd 147) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26349) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1908) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26219) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 10'sd 503) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11424) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13046) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19126) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14132) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3144) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14359) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1768) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28584) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4852) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18095) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11240) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2468) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26754) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4911) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_24[7:0]) +
	( 9'sd 148) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14471) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3783) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9328) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9163) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25707) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9769) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22889) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6975) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27904) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18500) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24529) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18038) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7841) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27562) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26821) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20420) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2757) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5278) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21172) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23080) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4232) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29271) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25751) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32720) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15568) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28166) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4818) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26454) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28146) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16558) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27191) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5887) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_78[7:0]) +
	( 10'sd 321) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24947) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20253) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22310) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_84[7:0]) +
	( 11'sd 678) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29150) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9711) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11106) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8471) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29362) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19483) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7864) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5399) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14900) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19058) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10559) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_102[7:0]) +
	( 12'sd 2014) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11077) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17473) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4692) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10882) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18729) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12147) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26585) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14094) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27613) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27573) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16780) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_122[7:0]) +
	( 11'sd 679) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6396) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11682) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22669) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 14'sd 6347) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31164) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7631) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23154) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31251) * $signed(input_fmap_5[7:0]) +
	( 11'sd 532) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12854) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20710) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20102) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24937) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22972) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15373) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6334) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10646) * $signed(input_fmap_16[7:0]) +
	( 10'sd 276) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28123) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_19[7:0]) +
	( 11'sd 633) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29354) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17031) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17743) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11709) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29068) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6029) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27446) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31462) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3136) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16279) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15648) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18277) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12399) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23654) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22957) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23263) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6956) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1530) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10113) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20371) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1990) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4700) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_52[7:0]) +
	( 11'sd 848) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15858) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17702) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25168) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9943) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1475) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12005) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26862) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24979) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25691) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1879) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24703) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16189) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24977) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19253) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18119) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3676) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3734) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16073) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24832) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8647) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31037) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19539) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3756) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20567) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1057) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29209) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13530) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30812) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32724) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21697) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5139) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15321) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31636) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32173) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20712) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10859) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10051) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 16'sd 25812) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11389) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13666) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10188) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24389) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7433) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2762) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22552) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9761) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26786) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1416) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10814) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16829) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30448) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29851) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25362) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16410) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29076) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30383) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_22[7:0]) +
	( 11'sd 578) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32240) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7698) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28950) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2426) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29127) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7614) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17878) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7240) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15978) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27410) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18948) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4476) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31941) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17383) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20833) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3364) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26063) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_54[7:0]) +
	( 11'sd 874) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9474) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25243) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29313) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26836) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25617) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1069) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20460) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4991) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16966) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32073) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14212) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19079) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31622) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11616) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23414) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31115) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14821) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28842) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30209) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11915) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14116) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13921) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21970) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_98[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17946) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20806) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21018) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20274) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25583) * $signed(input_fmap_105[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10079) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2153) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5346) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24887) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19495) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21137) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7113) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24530) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13953) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28793) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3695) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24926) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1303) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5793) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 16'sd 26362) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14186) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27784) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3125) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31186) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22437) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26821) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17075) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25675) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23213) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26647) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4599) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19823) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15994) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30053) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1701) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23510) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30602) * $signed(input_fmap_26[7:0]) +
	( 9'sd 130) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30757) * $signed(input_fmap_28[7:0]) +
	( 11'sd 745) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30550) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8787) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15649) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23062) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5120) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21774) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14650) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26320) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3663) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1662) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19765) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31178) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18920) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23760) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7395) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9578) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30493) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13292) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5346) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15449) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14744) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8194) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16165) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24858) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9753) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22744) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14171) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16160) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2458) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2737) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6255) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21473) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26233) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19074) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3256) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14734) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18736) * $signed(input_fmap_95[7:0]) +
	( 8'sd 105) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17090) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_98[7:0]) +
	( 11'sd 513) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7247) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23748) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31790) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24282) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24637) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23215) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_109[7:0]) +
	( 11'sd 972) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13449) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16432) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29699) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2975) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12341) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29045) * $signed(input_fmap_120[7:0]) +
	( 11'sd 672) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4388) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1518) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7213) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27556) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1542) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 16'sd 31907) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2840) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16938) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21140) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25894) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32024) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5342) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30140) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4708) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_14[7:0]) +
	( 11'sd 698) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8045) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32710) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19769) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10996) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30194) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27799) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26072) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23828) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30613) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15916) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15413) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1169) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21645) * $signed(input_fmap_42[7:0]) +
	( 11'sd 532) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22321) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23576) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27243) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1736) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29794) * $signed(input_fmap_55[7:0]) +
	( 6'sd 28) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18980) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19232) * $signed(input_fmap_59[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32615) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5354) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22110) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11304) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14017) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4125) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31744) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11069) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4715) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1824) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16781) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30176) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28493) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10912) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6611) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13607) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9533) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28947) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12702) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3101) * $signed(input_fmap_91[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18746) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18342) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22113) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14189) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12770) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30975) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20055) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18307) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12203) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10948) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7740) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1509) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12136) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16928) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25589) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19368) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26191) * $signed(input_fmap_114[7:0]) +
	( 6'sd 18) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9451) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16576) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14496) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2663) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3999) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26911) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14625) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30685) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 14'sd 4802) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8837) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_2[7:0]) +
	( 11'sd 784) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20536) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21145) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8350) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1411) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14986) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16051) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13455) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13972) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20918) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4658) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31562) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10325) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16627) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10125) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14692) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6421) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1352) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13751) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10036) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27011) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2108) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17485) * $signed(input_fmap_31[7:0]) +
	( 6'sd 19) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19980) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27546) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1674) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19883) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2674) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19875) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17920) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32242) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7424) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5867) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21404) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20263) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29976) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6454) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3173) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13620) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8926) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12677) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12281) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14367) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8607) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21342) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9872) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8328) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28219) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4733) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2301) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24221) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11871) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23571) * $signed(input_fmap_78[7:0]) +
	( 10'sd 287) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14877) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29332) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2212) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26917) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17622) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22208) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26093) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27370) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23274) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22902) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3801) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32218) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11802) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25692) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3479) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17074) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31801) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16616) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15434) * $signed(input_fmap_116[7:0]) +
	( 10'sd 322) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21842) * $signed(input_fmap_118[7:0]) +
	( 7'sd 55) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24204) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2468) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20738) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18931) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_125[7:0]) +
	( 12'sd 2027) * $signed(input_fmap_126[7:0]) +
	( 8'sd 82) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 16'sd 27681) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17036) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22283) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4599) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30594) * $signed(input_fmap_7[7:0]) +
	( 11'sd 613) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17273) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22678) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13067) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25219) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20748) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15358) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32204) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17826) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5729) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5186) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18501) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5071) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11290) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17963) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14963) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31172) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6979) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20529) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22277) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7722) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22002) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18379) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26642) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20786) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32105) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17175) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3441) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21342) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10335) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16234) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12704) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23521) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23518) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8484) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24066) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16136) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18907) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4330) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5966) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2933) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18352) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5635) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17116) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28053) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18714) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12979) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1909) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7231) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11104) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16828) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26211) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4390) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_86[7:0]) +
	( 11'sd 563) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20745) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15779) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9598) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1939) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12815) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2182) * $signed(input_fmap_96[7:0]) +
	( 10'sd 389) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1860) * $signed(input_fmap_98[7:0]) +
	( 11'sd 820) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24792) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3878) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8709) * $signed(input_fmap_103[7:0]) +
	( 10'sd 393) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14104) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23421) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7396) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20603) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30988) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_113[7:0]) +
	( 11'sd 576) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18429) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27577) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23827) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19351) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8244) * $signed(input_fmap_120[7:0]) +
	( 11'sd 551) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10561) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15302) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27086) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12669) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22460) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 15'sd 9054) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29673) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2578) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18155) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_7[7:0]) +
	( 11'sd 534) * $signed(input_fmap_8[7:0]) +
	( 10'sd 279) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8404) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18904) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10204) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12789) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12469) * $signed(input_fmap_16[7:0]) +
	( 10'sd 317) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8524) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32613) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5524) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26638) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7022) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1335) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6098) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17394) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21530) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32282) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14311) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14307) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2805) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3448) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32534) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28763) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5574) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12304) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24650) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29640) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16780) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7606) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29571) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25163) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3863) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23282) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32619) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24705) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7721) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_66[7:0]) +
	( 13'sd 4003) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10406) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5131) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1401) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23620) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14130) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24400) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18533) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31108) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7640) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10104) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7100) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18918) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16817) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1411) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9072) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28310) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17701) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4193) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28871) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18392) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23877) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17518) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13111) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18420) * $signed(input_fmap_101[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8830) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28901) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27622) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10449) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27539) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25097) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18155) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_113[7:0]) +
	( 11'sd 902) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22524) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7844) * $signed(input_fmap_117[7:0]) +
	( 14'sd 8092) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8301) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15068) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26852) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21460) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1377) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9139) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19139) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13798) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 14'sd 7658) * $signed(input_fmap_0[7:0]) +
	( 10'sd 505) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15028) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7116) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28534) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5032) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10749) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14970) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7868) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28264) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31508) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12569) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25917) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7073) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1574) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1211) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1456) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11949) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19038) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21114) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28612) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8939) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31745) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13467) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28614) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16236) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23916) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11732) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12833) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5581) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8809) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28241) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16974) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25972) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17076) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22371) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12399) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25940) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1609) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10867) * $signed(input_fmap_67[7:0]) +
	( 10'sd 470) * $signed(input_fmap_68[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20059) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26165) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26707) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16912) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27187) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20615) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28144) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27250) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30922) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10569) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20751) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22092) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_89[7:0]) +
	( 10'sd 400) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11392) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29536) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_99[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10716) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30407) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_104[7:0]) +
	( 11'sd 687) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_106[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10145) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_110[7:0]) +
	( 8'sd 101) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28585) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28328) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13530) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18252) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25903) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11856) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23273) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13068) * $signed(input_fmap_123[7:0]) +
	( 10'sd 291) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6208) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_126[7:0]) +
	( 11'sd 560) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 16'sd 32327) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13309) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11387) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8694) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20735) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10794) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26114) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7347) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31511) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6175) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4356) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13052) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5535) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_21[7:0]) +
	( 10'sd 332) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9090) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27222) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27101) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31714) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23285) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12129) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31704) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4227) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15002) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4219) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17973) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22519) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16816) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21832) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6407) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31298) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2322) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31652) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9215) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20361) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32639) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4521) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30781) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1765) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32543) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20257) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2445) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20844) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26882) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24616) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24973) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15548) * $signed(input_fmap_68[7:0]) +
	( 10'sd 404) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15088) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29938) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29302) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11106) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5344) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2643) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7899) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30948) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15693) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27784) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8829) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13981) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9439) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29751) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29817) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32708) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21910) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29795) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23865) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19701) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8376) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4751) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2057) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25124) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25206) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20173) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5672) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24592) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22549) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3709) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25351) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17998) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10189) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29663) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20327) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6568) * $signed(input_fmap_124[7:0]) +
	( 9'sd 187) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 15'sd 10909) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27304) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2145) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26602) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16754) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4292) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3274) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5570) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27972) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7778) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13149) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5672) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15313) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7983) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11984) * $signed(input_fmap_23[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17307) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25153) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20417) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5645) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1271) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11308) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27402) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10072) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23102) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24087) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10951) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14075) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18633) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11334) * $signed(input_fmap_47[7:0]) +
	( 11'sd 610) * $signed(input_fmap_48[7:0]) +
	( 11'sd 895) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32595) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19147) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3482) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29148) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14609) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28213) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31397) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_60[7:0]) +
	( 11'sd 526) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11412) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16690) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30500) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19504) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24452) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19644) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17145) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9584) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10518) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17439) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15834) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12730) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6532) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24709) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3669) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17926) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22209) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3672) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18863) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27853) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16121) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5825) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31628) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29627) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31455) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10919) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12760) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26280) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_106[7:0]) +
	( 9'sd 189) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7983) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24548) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20177) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8598) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11807) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18696) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7253) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21139) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27739) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31985) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15291) * $signed(input_fmap_123[7:0]) +
	( 7'sd 32) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23237) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31773) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23757) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 13'sd 2452) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20019) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22126) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4225) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32114) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9088) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5576) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14421) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16872) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9095) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21311) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10300) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4104) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11238) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23462) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2884) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4734) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25763) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26921) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20136) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3683) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4370) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13760) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12449) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21437) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21597) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24306) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2833) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_50[7:0]) +
	( 9'sd 219) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17757) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17988) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7032) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20660) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24141) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16424) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13687) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22048) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15203) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13462) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28916) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10049) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16983) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30756) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20595) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15188) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2920) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15921) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27155) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21289) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13387) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23474) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11734) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24379) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16528) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27891) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2996) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17635) * $signed(input_fmap_87[7:0]) +
	( 11'sd 993) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16007) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_91[7:0]) +
	( 11'sd 532) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32220) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23865) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2348) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27072) * $signed(input_fmap_100[7:0]) +
	( 8'sd 64) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30078) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28923) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28606) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28002) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18612) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31532) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24202) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9773) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5773) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2166) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6568) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21300) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13476) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16582) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18672) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13715) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9499) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31756) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 16'sd 26170) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2728) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8185) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30765) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22335) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21138) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22376) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10946) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14225) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11957) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11805) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30064) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5378) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23553) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30152) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3960) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23123) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25306) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7302) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25112) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21084) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28372) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30823) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8320) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26446) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29027) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2182) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21791) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5682) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18843) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24659) * $signed(input_fmap_48[7:0]) +
	( 11'sd 976) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30032) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12310) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17261) * $signed(input_fmap_52[7:0]) +
	( 10'sd 379) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_54[7:0]) +
	( 12'sd 2033) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5946) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4276) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18863) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15525) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13483) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2523) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23335) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32636) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32113) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4755) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1045) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10346) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23967) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25160) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3009) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10829) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21928) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16007) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25655) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28904) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16198) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5609) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16782) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15839) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30510) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12912) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17798) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31623) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3643) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24225) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27277) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24870) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9214) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15304) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21207) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26426) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31600) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19352) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9304) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7909) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15059) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20887) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1319) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10337) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_127[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 16'd20052;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 16'd23139;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 16'd20912;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 15'd14176;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 15'd8354;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 15'd11449;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 12'd1076;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 16'd27718;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 16'd29878;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 15'd15765;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 14'd5953;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 16'd22409;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 16'd20652;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 16'd23506;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 16'd21989;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 16'd27744;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 14'd7482;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 16'd18529;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 14'd5718;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 15'd11425;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 15'd14173;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 16'd22089;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 15'd14422;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 12'd2042;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 15'd8368;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 16'd19686;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 16'd29138;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 16'd28437;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 12'd1184;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 11'd615;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 16'd16483;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 11'd893;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 14'd7702;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 16'd23856;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 14'd6171;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 16'd19713;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 15'd16222;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 15'd14468;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 16'd18421;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 14'd6644;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 15'd15699;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 15'd8844;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 14'd4185;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 16'd22658;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 16'd20469;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 16'd19680;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 14'd8011;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 15'd13777;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 16'd32361;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 16'd30142;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 16'd22217;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 16'd20111;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 15'd12871;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 13'd2389;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 16'd29170;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 16'd26117;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 10'd323;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 14'd6648;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 16'd17245;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 16'd18061;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 13'd3944;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 16'd30129;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 14'd7935;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 14'd5199;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 13'd2462;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 15'd10150;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 16'd25345;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 15'd10195;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 11'd587;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 11'd702;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 14'd4953;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 16'd23149;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 16'd32164;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 15'd15627;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 15'd8527;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 16'd29327;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 13'd2071;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 15'd13213;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 15'd13966;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 16'd31368;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 16'd30282;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 16'd16577;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 16'd32048;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 15'd14002;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 16'd23126;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 15'd9328;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 14'd6888;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 16'd17334;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 16'd26919;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 16'd17345;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 16'd19288;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 15'd12904;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 16'd17998;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 15'd11056;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 15'd9833;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 15'd12439;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 16'd26075;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 16'd26537;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 16'd32235;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 16'd27441;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 16'd23166;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 16'd17465;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 9'd245;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 15'd10791;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 16'd28484;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 14'd6003;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 16'd29893;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 16'd22743;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 16'd23700;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 12'd1976;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 16'd23913;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 15'd13235;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 16'd25354;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 16'd19159;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 15'd9012;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 13'd3104;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 16'd28744;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 16'd18948;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 15'd11943;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 16'd25389;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 16'd20375;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 16'd21465;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 15'd13251;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 16'd31307;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 16'd31884;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 16'd30154;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 15'd12121;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 14'd6697;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[21:15]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[21:15]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[21:15]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[21:15]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[21:15]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[21:15]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[21:15]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[21:15]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[21:15]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[21:15]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[21:15]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[21:15]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[21:15]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[21:15]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[21:15]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[21:15]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[21:15]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[21:15]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[21:15]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[21:15]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[21:15]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[21:15]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[21:15]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[21:15]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[21:15]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[21:15]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[21:15]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[21:15]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[21:15]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[21:15]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[21:15]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[21:15]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[21:15]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[21:15]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[21:15]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[21:15]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[21:15]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[21:15]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[21:15]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[21:15]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[21:15]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[21:15]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[21:15]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[21:15]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[21:15]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[21:15]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[21:15]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[21:15]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[21:15]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[21:15]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[21:15]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[21:15]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[21:15]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[21:15]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[21:15]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[21:15]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[21:15]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[21:15]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[21:15]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[21:15]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[21:15]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[21:15]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[21:15]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[21:15]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[21:15]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[21:15]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[21:15]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[21:15]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[21:15]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[21:15]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[21:15]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[21:15]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[21:15]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[21:15]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[21:15]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[21:15]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[21:15]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[21:15]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[21:15]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[21:15]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[21:15]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[21:15]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[21:15]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[21:15]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[21:15]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[21:15]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[21:15]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[21:15]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[21:15]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[21:15]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[21:15]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[21:15]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[21:15]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[21:15]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[21:15]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[21:15]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[21:15]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[21:15]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[21:15]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[21:15]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[21:15]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[21:15]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[21:15]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[21:15]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[21:15]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[21:15]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[21:15]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[21:15]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[21:15]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[21:15]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[21:15]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[21:15]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[21:15]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[21:15]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[21:15]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[21:15]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[21:15]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[21:15]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[21:15]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[21:15]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[21:15]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[21:15]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[21:15]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[21:15]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[21:15]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[21:15]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[21:15]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[21:15]}} :'d6) : '0;

assign output_act = {
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
