module conv14_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [2048-1:0] input_act,
    output logic [2048-1:0] output_act,
    output logic ready
);

logic [2048-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];
logic [7:0] input_fmap_128;
assign input_fmap_128 = input_act_ff[1031:1024];
logic [7:0] input_fmap_129;
assign input_fmap_129 = input_act_ff[1039:1032];
logic [7:0] input_fmap_130;
assign input_fmap_130 = input_act_ff[1047:1040];
logic [7:0] input_fmap_131;
assign input_fmap_131 = input_act_ff[1055:1048];
logic [7:0] input_fmap_132;
assign input_fmap_132 = input_act_ff[1063:1056];
logic [7:0] input_fmap_133;
assign input_fmap_133 = input_act_ff[1071:1064];
logic [7:0] input_fmap_134;
assign input_fmap_134 = input_act_ff[1079:1072];
logic [7:0] input_fmap_135;
assign input_fmap_135 = input_act_ff[1087:1080];
logic [7:0] input_fmap_136;
assign input_fmap_136 = input_act_ff[1095:1088];
logic [7:0] input_fmap_137;
assign input_fmap_137 = input_act_ff[1103:1096];
logic [7:0] input_fmap_138;
assign input_fmap_138 = input_act_ff[1111:1104];
logic [7:0] input_fmap_139;
assign input_fmap_139 = input_act_ff[1119:1112];
logic [7:0] input_fmap_140;
assign input_fmap_140 = input_act_ff[1127:1120];
logic [7:0] input_fmap_141;
assign input_fmap_141 = input_act_ff[1135:1128];
logic [7:0] input_fmap_142;
assign input_fmap_142 = input_act_ff[1143:1136];
logic [7:0] input_fmap_143;
assign input_fmap_143 = input_act_ff[1151:1144];
logic [7:0] input_fmap_144;
assign input_fmap_144 = input_act_ff[1159:1152];
logic [7:0] input_fmap_145;
assign input_fmap_145 = input_act_ff[1167:1160];
logic [7:0] input_fmap_146;
assign input_fmap_146 = input_act_ff[1175:1168];
logic [7:0] input_fmap_147;
assign input_fmap_147 = input_act_ff[1183:1176];
logic [7:0] input_fmap_148;
assign input_fmap_148 = input_act_ff[1191:1184];
logic [7:0] input_fmap_149;
assign input_fmap_149 = input_act_ff[1199:1192];
logic [7:0] input_fmap_150;
assign input_fmap_150 = input_act_ff[1207:1200];
logic [7:0] input_fmap_151;
assign input_fmap_151 = input_act_ff[1215:1208];
logic [7:0] input_fmap_152;
assign input_fmap_152 = input_act_ff[1223:1216];
logic [7:0] input_fmap_153;
assign input_fmap_153 = input_act_ff[1231:1224];
logic [7:0] input_fmap_154;
assign input_fmap_154 = input_act_ff[1239:1232];
logic [7:0] input_fmap_155;
assign input_fmap_155 = input_act_ff[1247:1240];
logic [7:0] input_fmap_156;
assign input_fmap_156 = input_act_ff[1255:1248];
logic [7:0] input_fmap_157;
assign input_fmap_157 = input_act_ff[1263:1256];
logic [7:0] input_fmap_158;
assign input_fmap_158 = input_act_ff[1271:1264];
logic [7:0] input_fmap_159;
assign input_fmap_159 = input_act_ff[1279:1272];
logic [7:0] input_fmap_160;
assign input_fmap_160 = input_act_ff[1287:1280];
logic [7:0] input_fmap_161;
assign input_fmap_161 = input_act_ff[1295:1288];
logic [7:0] input_fmap_162;
assign input_fmap_162 = input_act_ff[1303:1296];
logic [7:0] input_fmap_163;
assign input_fmap_163 = input_act_ff[1311:1304];
logic [7:0] input_fmap_164;
assign input_fmap_164 = input_act_ff[1319:1312];
logic [7:0] input_fmap_165;
assign input_fmap_165 = input_act_ff[1327:1320];
logic [7:0] input_fmap_166;
assign input_fmap_166 = input_act_ff[1335:1328];
logic [7:0] input_fmap_167;
assign input_fmap_167 = input_act_ff[1343:1336];
logic [7:0] input_fmap_168;
assign input_fmap_168 = input_act_ff[1351:1344];
logic [7:0] input_fmap_169;
assign input_fmap_169 = input_act_ff[1359:1352];
logic [7:0] input_fmap_170;
assign input_fmap_170 = input_act_ff[1367:1360];
logic [7:0] input_fmap_171;
assign input_fmap_171 = input_act_ff[1375:1368];
logic [7:0] input_fmap_172;
assign input_fmap_172 = input_act_ff[1383:1376];
logic [7:0] input_fmap_173;
assign input_fmap_173 = input_act_ff[1391:1384];
logic [7:0] input_fmap_174;
assign input_fmap_174 = input_act_ff[1399:1392];
logic [7:0] input_fmap_175;
assign input_fmap_175 = input_act_ff[1407:1400];
logic [7:0] input_fmap_176;
assign input_fmap_176 = input_act_ff[1415:1408];
logic [7:0] input_fmap_177;
assign input_fmap_177 = input_act_ff[1423:1416];
logic [7:0] input_fmap_178;
assign input_fmap_178 = input_act_ff[1431:1424];
logic [7:0] input_fmap_179;
assign input_fmap_179 = input_act_ff[1439:1432];
logic [7:0] input_fmap_180;
assign input_fmap_180 = input_act_ff[1447:1440];
logic [7:0] input_fmap_181;
assign input_fmap_181 = input_act_ff[1455:1448];
logic [7:0] input_fmap_182;
assign input_fmap_182 = input_act_ff[1463:1456];
logic [7:0] input_fmap_183;
assign input_fmap_183 = input_act_ff[1471:1464];
logic [7:0] input_fmap_184;
assign input_fmap_184 = input_act_ff[1479:1472];
logic [7:0] input_fmap_185;
assign input_fmap_185 = input_act_ff[1487:1480];
logic [7:0] input_fmap_186;
assign input_fmap_186 = input_act_ff[1495:1488];
logic [7:0] input_fmap_187;
assign input_fmap_187 = input_act_ff[1503:1496];
logic [7:0] input_fmap_188;
assign input_fmap_188 = input_act_ff[1511:1504];
logic [7:0] input_fmap_189;
assign input_fmap_189 = input_act_ff[1519:1512];
logic [7:0] input_fmap_190;
assign input_fmap_190 = input_act_ff[1527:1520];
logic [7:0] input_fmap_191;
assign input_fmap_191 = input_act_ff[1535:1528];
logic [7:0] input_fmap_192;
assign input_fmap_192 = input_act_ff[1543:1536];
logic [7:0] input_fmap_193;
assign input_fmap_193 = input_act_ff[1551:1544];
logic [7:0] input_fmap_194;
assign input_fmap_194 = input_act_ff[1559:1552];
logic [7:0] input_fmap_195;
assign input_fmap_195 = input_act_ff[1567:1560];
logic [7:0] input_fmap_196;
assign input_fmap_196 = input_act_ff[1575:1568];
logic [7:0] input_fmap_197;
assign input_fmap_197 = input_act_ff[1583:1576];
logic [7:0] input_fmap_198;
assign input_fmap_198 = input_act_ff[1591:1584];
logic [7:0] input_fmap_199;
assign input_fmap_199 = input_act_ff[1599:1592];
logic [7:0] input_fmap_200;
assign input_fmap_200 = input_act_ff[1607:1600];
logic [7:0] input_fmap_201;
assign input_fmap_201 = input_act_ff[1615:1608];
logic [7:0] input_fmap_202;
assign input_fmap_202 = input_act_ff[1623:1616];
logic [7:0] input_fmap_203;
assign input_fmap_203 = input_act_ff[1631:1624];
logic [7:0] input_fmap_204;
assign input_fmap_204 = input_act_ff[1639:1632];
logic [7:0] input_fmap_205;
assign input_fmap_205 = input_act_ff[1647:1640];
logic [7:0] input_fmap_206;
assign input_fmap_206 = input_act_ff[1655:1648];
logic [7:0] input_fmap_207;
assign input_fmap_207 = input_act_ff[1663:1656];
logic [7:0] input_fmap_208;
assign input_fmap_208 = input_act_ff[1671:1664];
logic [7:0] input_fmap_209;
assign input_fmap_209 = input_act_ff[1679:1672];
logic [7:0] input_fmap_210;
assign input_fmap_210 = input_act_ff[1687:1680];
logic [7:0] input_fmap_211;
assign input_fmap_211 = input_act_ff[1695:1688];
logic [7:0] input_fmap_212;
assign input_fmap_212 = input_act_ff[1703:1696];
logic [7:0] input_fmap_213;
assign input_fmap_213 = input_act_ff[1711:1704];
logic [7:0] input_fmap_214;
assign input_fmap_214 = input_act_ff[1719:1712];
logic [7:0] input_fmap_215;
assign input_fmap_215 = input_act_ff[1727:1720];
logic [7:0] input_fmap_216;
assign input_fmap_216 = input_act_ff[1735:1728];
logic [7:0] input_fmap_217;
assign input_fmap_217 = input_act_ff[1743:1736];
logic [7:0] input_fmap_218;
assign input_fmap_218 = input_act_ff[1751:1744];
logic [7:0] input_fmap_219;
assign input_fmap_219 = input_act_ff[1759:1752];
logic [7:0] input_fmap_220;
assign input_fmap_220 = input_act_ff[1767:1760];
logic [7:0] input_fmap_221;
assign input_fmap_221 = input_act_ff[1775:1768];
logic [7:0] input_fmap_222;
assign input_fmap_222 = input_act_ff[1783:1776];
logic [7:0] input_fmap_223;
assign input_fmap_223 = input_act_ff[1791:1784];
logic [7:0] input_fmap_224;
assign input_fmap_224 = input_act_ff[1799:1792];
logic [7:0] input_fmap_225;
assign input_fmap_225 = input_act_ff[1807:1800];
logic [7:0] input_fmap_226;
assign input_fmap_226 = input_act_ff[1815:1808];
logic [7:0] input_fmap_227;
assign input_fmap_227 = input_act_ff[1823:1816];
logic [7:0] input_fmap_228;
assign input_fmap_228 = input_act_ff[1831:1824];
logic [7:0] input_fmap_229;
assign input_fmap_229 = input_act_ff[1839:1832];
logic [7:0] input_fmap_230;
assign input_fmap_230 = input_act_ff[1847:1840];
logic [7:0] input_fmap_231;
assign input_fmap_231 = input_act_ff[1855:1848];
logic [7:0] input_fmap_232;
assign input_fmap_232 = input_act_ff[1863:1856];
logic [7:0] input_fmap_233;
assign input_fmap_233 = input_act_ff[1871:1864];
logic [7:0] input_fmap_234;
assign input_fmap_234 = input_act_ff[1879:1872];
logic [7:0] input_fmap_235;
assign input_fmap_235 = input_act_ff[1887:1880];
logic [7:0] input_fmap_236;
assign input_fmap_236 = input_act_ff[1895:1888];
logic [7:0] input_fmap_237;
assign input_fmap_237 = input_act_ff[1903:1896];
logic [7:0] input_fmap_238;
assign input_fmap_238 = input_act_ff[1911:1904];
logic [7:0] input_fmap_239;
assign input_fmap_239 = input_act_ff[1919:1912];
logic [7:0] input_fmap_240;
assign input_fmap_240 = input_act_ff[1927:1920];
logic [7:0] input_fmap_241;
assign input_fmap_241 = input_act_ff[1935:1928];
logic [7:0] input_fmap_242;
assign input_fmap_242 = input_act_ff[1943:1936];
logic [7:0] input_fmap_243;
assign input_fmap_243 = input_act_ff[1951:1944];
logic [7:0] input_fmap_244;
assign input_fmap_244 = input_act_ff[1959:1952];
logic [7:0] input_fmap_245;
assign input_fmap_245 = input_act_ff[1967:1960];
logic [7:0] input_fmap_246;
assign input_fmap_246 = input_act_ff[1975:1968];
logic [7:0] input_fmap_247;
assign input_fmap_247 = input_act_ff[1983:1976];
logic [7:0] input_fmap_248;
assign input_fmap_248 = input_act_ff[1991:1984];
logic [7:0] input_fmap_249;
assign input_fmap_249 = input_act_ff[1999:1992];
logic [7:0] input_fmap_250;
assign input_fmap_250 = input_act_ff[2007:2000];
logic [7:0] input_fmap_251;
assign input_fmap_251 = input_act_ff[2015:2008];
logic [7:0] input_fmap_252;
assign input_fmap_252 = input_act_ff[2023:2016];
logic [7:0] input_fmap_253;
assign input_fmap_253 = input_act_ff[2031:2024];
logic [7:0] input_fmap_254;
assign input_fmap_254 = input_act_ff[2039:2032];
logic [7:0] input_fmap_255;
assign input_fmap_255 = input_act_ff[2047:2040];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_128;
assign conv_mac_128 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_129;
assign conv_mac_129 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_130;
assign conv_mac_130 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_131;
assign conv_mac_131 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_132;
assign conv_mac_132 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_133;
assign conv_mac_133 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_134;
assign conv_mac_134 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_135;
assign conv_mac_135 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_136;
assign conv_mac_136 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_137;
assign conv_mac_137 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_138;
assign conv_mac_138 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_139;
assign conv_mac_139 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_140;
assign conv_mac_140 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_141;
assign conv_mac_141 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_142;
assign conv_mac_142 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_143;
assign conv_mac_143 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_144;
assign conv_mac_144 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_145;
assign conv_mac_145 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_146;
assign conv_mac_146 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_147;
assign conv_mac_147 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_148;
assign conv_mac_148 = 
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_149;
assign conv_mac_149 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_150;
assign conv_mac_150 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_151;
assign conv_mac_151 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_152;
assign conv_mac_152 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_153;
assign conv_mac_153 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_154;
assign conv_mac_154 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_155;
assign conv_mac_155 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_156;
assign conv_mac_156 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_157;
assign conv_mac_157 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_158;
assign conv_mac_158 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_159;
assign conv_mac_159 = 
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_160;
assign conv_mac_160 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_161;
assign conv_mac_161 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_162;
assign conv_mac_162 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_163;
assign conv_mac_163 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_164;
assign conv_mac_164 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_165;
assign conv_mac_165 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_166;
assign conv_mac_166 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_167;
assign conv_mac_167 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_168;
assign conv_mac_168 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_169;
assign conv_mac_169 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_170;
assign conv_mac_170 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_171;
assign conv_mac_171 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_172;
assign conv_mac_172 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_173;
assign conv_mac_173 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_174;
assign conv_mac_174 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_175;
assign conv_mac_175 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_176;
assign conv_mac_176 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_177;
assign conv_mac_177 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_178;
assign conv_mac_178 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_179;
assign conv_mac_179 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_180;
assign conv_mac_180 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_181;
assign conv_mac_181 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_182;
assign conv_mac_182 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_183;
assign conv_mac_183 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_184;
assign conv_mac_184 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_185;
assign conv_mac_185 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_186;
assign conv_mac_186 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_187;
assign conv_mac_187 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_188;
assign conv_mac_188 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_189;
assign conv_mac_189 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_190;
assign conv_mac_190 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_191;
assign conv_mac_191 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_192;
assign conv_mac_192 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_193;
assign conv_mac_193 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_194;
assign conv_mac_194 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_195;
assign conv_mac_195 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_196;
assign conv_mac_196 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_197;
assign conv_mac_197 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_198;
assign conv_mac_198 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_199;
assign conv_mac_199 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_200;
assign conv_mac_200 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_201;
assign conv_mac_201 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_202;
assign conv_mac_202 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_203;
assign conv_mac_203 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_204;
assign conv_mac_204 = 
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_205;
assign conv_mac_205 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_206;
assign conv_mac_206 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_207;
assign conv_mac_207 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_208;
assign conv_mac_208 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]);

logic signed [31:0] conv_mac_209;
assign conv_mac_209 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]);

logic signed [31:0] conv_mac_210;
assign conv_mac_210 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_211;
assign conv_mac_211 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_212;
assign conv_mac_212 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_213;
assign conv_mac_213 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_214;
assign conv_mac_214 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_215;
assign conv_mac_215 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_216;
assign conv_mac_216 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_217;
assign conv_mac_217 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_218;
assign conv_mac_218 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_219;
assign conv_mac_219 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_220;
assign conv_mac_220 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_221;
assign conv_mac_221 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_222;
assign conv_mac_222 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_223;
assign conv_mac_223 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_224;
assign conv_mac_224 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_225;
assign conv_mac_225 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_226;
assign conv_mac_226 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_227;
assign conv_mac_227 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_228;
assign conv_mac_228 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_229;
assign conv_mac_229 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_230;
assign conv_mac_230 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_231;
assign conv_mac_231 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_232;
assign conv_mac_232 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_233;
assign conv_mac_233 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_234;
assign conv_mac_234 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_235;
assign conv_mac_235 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_236;
assign conv_mac_236 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_237;
assign conv_mac_237 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_238;
assign conv_mac_238 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 3'sd 2) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_239;
assign conv_mac_239 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_240;
assign conv_mac_240 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_241;
assign conv_mac_241 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_242;
assign conv_mac_242 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_243;
assign conv_mac_243 = 
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 3'sd 2) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_244;
assign conv_mac_244 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 3'sd 2) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_194[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_245;
assign conv_mac_245 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 3'sd 2) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 3'sd 2) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]);

logic signed [31:0] conv_mac_246;
assign conv_mac_246 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 3'sd 2) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 3'sd 2) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_247;
assign conv_mac_247 = 
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 3'sd 2) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 3'sd 2) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 3'sd 2) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 3'sd 2) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_248;
assign conv_mac_248 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_150[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 3'sd 2) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 3'sd 2) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 3'sd 2) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_249;
assign conv_mac_249 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 3'sd 2) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 3'sd 2) * $signed(input_fmap_174[7:0]) +
	( 3'sd 2) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 3'sd 2) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_250;
assign conv_mac_250 = 
	( 3'sd 2) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 3'sd 2) * $signed(input_fmap_16[7:0]) +
	( 3'sd 2) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 3'sd 2) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 3'sd 2) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_36[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 3'sd 2) * $signed(input_fmap_47[7:0]) +
	( 3'sd 2) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 3'sd 2) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_65[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 3'sd 2) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 3'sd 2) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 3'sd 2) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 3'sd 2) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 3'sd 2) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 3'sd 2) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_251;
assign conv_mac_251 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_9[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 3'sd 2) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 3'sd 2) * $signed(input_fmap_25[7:0]) +
	( 3'sd 2) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 3'sd 2) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 3'sd 2) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 3'sd 2) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 2'sd 1) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 3'sd 2) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 2'sd 1) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 2'sd 1) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 3'sd 2) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_115[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 2'sd 1) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 3'sd 2) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_194[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 3'sd 2) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 3'sd 2) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 3'sd 2) * $signed(input_fmap_227[7:0]) +
	( 3'sd 2) * $signed(input_fmap_228[7:0]) +
	( 3'sd 2) * $signed(input_fmap_229[7:0]) +
	( 3'sd 2) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_252;
assign conv_mac_252 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 2'sd 1) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 3'sd 2) * $signed(input_fmap_30[7:0]) +
	( 3'sd 2) * $signed(input_fmap_33[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 3'sd 2) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 3'sd 2) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_60[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 3'sd 2) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_65[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 3'sd 2) * $signed(input_fmap_71[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 3'sd 2) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_89[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_92[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 3'sd 2) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_115[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 3'sd 2) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 3'sd 2) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 2'sd 1) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 2'sd 1) * $signed(input_fmap_168[7:0]) +
	( 2'sd 1) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 2'sd 1) * $signed(input_fmap_184[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 3'sd 2) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 2'sd 1) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_213[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 3'sd 2) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_253;
assign conv_mac_253 = 
	( 2'sd 1) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 3'sd 2) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_9[7:0]) +
	( 3'sd 2) * $signed(input_fmap_10[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_15[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_18[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_34[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 2'sd 1) * $signed(input_fmap_36[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 3'sd 2) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 3'sd 2) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 3'sd 2) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_61[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 3'sd 2) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 2'sd 1) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 2'sd 1) * $signed(input_fmap_88[7:0]) +
	( 2'sd 1) * $signed(input_fmap_90[7:0]) +
	( 2'sd 1) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 3'sd 2) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 3'sd 2) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 3'sd 2) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 2'sd 1) * $signed(input_fmap_107[7:0]) +
	( 3'sd 2) * $signed(input_fmap_108[7:0]) +
	( 3'sd 2) * $signed(input_fmap_109[7:0]) +
	( 3'sd 2) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_112[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 3'sd 2) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 3'sd 2) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_141[7:0]) +
	( 3'sd 2) * $signed(input_fmap_142[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_146[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 2'sd 1) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 2'sd 1) * $signed(input_fmap_150[7:0]) +
	( 2'sd 1) * $signed(input_fmap_151[7:0]) +
	( 2'sd 1) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 2'sd 1) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_159[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_170[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 3'sd 2) * $signed(input_fmap_177[7:0]) +
	( 3'sd 2) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_190[7:0]) +
	( 3'sd 2) * $signed(input_fmap_191[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_198[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 3'sd 2) * $signed(input_fmap_200[7:0]) +
	( 3'sd 2) * $signed(input_fmap_201[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 3'sd 2) * $signed(input_fmap_204[7:0]) +
	( 3'sd 2) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 2'sd 1) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_224[7:0]) +
	( 3'sd 2) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_227[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 3'sd 2) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_233[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_236[7:0]) +
	( 3'sd 2) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 3'sd 2) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_240[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 3'sd 2) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 2'sd 1) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_251[7:0]) +
	( 2'sd 1) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 2'sd 1) * $signed(input_fmap_254[7:0]) +
	( 3'sd 2) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_254;
assign conv_mac_254 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 3'sd 2) * $signed(input_fmap_3[7:0]) +
	( 3'sd 2) * $signed(input_fmap_4[7:0]) +
	( 2'sd 1) * $signed(input_fmap_5[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 2'sd 1) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 3'sd 2) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_13[7:0]) +
	( 3'sd 2) * $signed(input_fmap_14[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 2'sd 1) * $signed(input_fmap_19[7:0]) +
	( 2'sd 1) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_21[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 3'sd 2) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 3'sd 2) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_30[7:0]) +
	( 2'sd 1) * $signed(input_fmap_33[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 3'sd 2) * $signed(input_fmap_38[7:0]) +
	( 3'sd 2) * $signed(input_fmap_39[7:0]) +
	( 3'sd 2) * $signed(input_fmap_40[7:0]) +
	( 2'sd 1) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_46[7:0]) +
	( 2'sd 1) * $signed(input_fmap_47[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_49[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_52[7:0]) +
	( 2'sd 1) * $signed(input_fmap_53[7:0]) +
	( 3'sd 2) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_55[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 3'sd 2) * $signed(input_fmap_61[7:0]) +
	( 3'sd 2) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 2'sd 1) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_68[7:0]) +
	( 3'sd 2) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 3'sd 2) * $signed(input_fmap_72[7:0]) +
	( 3'sd 2) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 2'sd 1) * $signed(input_fmap_78[7:0]) +
	( 3'sd 2) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 3'sd 2) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_88[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 2'sd 1) * $signed(input_fmap_93[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 2'sd 1) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_108[7:0]) +
	( 2'sd 1) * $signed(input_fmap_109[7:0]) +
	( 2'sd 1) * $signed(input_fmap_110[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 2'sd 1) * $signed(input_fmap_113[7:0]) +
	( 2'sd 1) * $signed(input_fmap_114[7:0]) +
	( 2'sd 1) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 2'sd 1) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 3'sd 2) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_127[7:0]) +
	( 3'sd 2) * $signed(input_fmap_128[7:0]) +
	( 2'sd 1) * $signed(input_fmap_129[7:0]) +
	( 2'sd 1) * $signed(input_fmap_130[7:0]) +
	( 3'sd 2) * $signed(input_fmap_131[7:0]) +
	( 2'sd 1) * $signed(input_fmap_132[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 3'sd 2) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_136[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 3'sd 2) * $signed(input_fmap_140[7:0]) +
	( 2'sd 1) * $signed(input_fmap_143[7:0]) +
	( 2'sd 1) * $signed(input_fmap_144[7:0]) +
	( 2'sd 1) * $signed(input_fmap_145[7:0]) +
	( 3'sd 2) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_148[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_159[7:0]) +
	( 2'sd 1) * $signed(input_fmap_160[7:0]) +
	( 3'sd 2) * $signed(input_fmap_161[7:0]) +
	( 3'sd 2) * $signed(input_fmap_162[7:0]) +
	( 2'sd 1) * $signed(input_fmap_163[7:0]) +
	( 2'sd 1) * $signed(input_fmap_164[7:0]) +
	( 3'sd 2) * $signed(input_fmap_165[7:0]) +
	( 2'sd 1) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 3'sd 2) * $signed(input_fmap_170[7:0]) +
	( 3'sd 2) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 3'sd 2) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_174[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 3'sd 2) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 3'sd 2) * $signed(input_fmap_182[7:0]) +
	( 3'sd 2) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_184[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_187[7:0]) +
	( 3'sd 2) * $signed(input_fmap_188[7:0]) +
	( 2'sd 1) * $signed(input_fmap_189[7:0]) +
	( 3'sd 2) * $signed(input_fmap_190[7:0]) +
	( 2'sd 1) * $signed(input_fmap_191[7:0]) +
	( 3'sd 2) * $signed(input_fmap_192[7:0]) +
	( 2'sd 1) * $signed(input_fmap_193[7:0]) +
	( 3'sd 2) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 3'sd 2) * $signed(input_fmap_197[7:0]) +
	( 2'sd 1) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_201[7:0]) +
	( 3'sd 2) * $signed(input_fmap_202[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 2'sd 1) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_209[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_213[7:0]) +
	( 2'sd 1) * $signed(input_fmap_214[7:0]) +
	( 3'sd 2) * $signed(input_fmap_215[7:0]) +
	( 2'sd 1) * $signed(input_fmap_216[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_218[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_220[7:0]) +
	( 3'sd 2) * $signed(input_fmap_221[7:0]) +
	( 2'sd 1) * $signed(input_fmap_222[7:0]) +
	( 3'sd 2) * $signed(input_fmap_224[7:0]) +
	( 2'sd 1) * $signed(input_fmap_226[7:0]) +
	( 2'sd 1) * $signed(input_fmap_228[7:0]) +
	( 2'sd 1) * $signed(input_fmap_229[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 3'sd 2) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 2'sd 1) * $signed(input_fmap_235[7:0]) +
	( 3'sd 2) * $signed(input_fmap_236[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 3'sd 2) * $signed(input_fmap_242[7:0]) +
	( 3'sd 2) * $signed(input_fmap_243[7:0]) +
	( 2'sd 1) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 3'sd 2) * $signed(input_fmap_248[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 2'sd 1) * $signed(input_fmap_253[7:0]) +
	( 3'sd 2) * $signed(input_fmap_254[7:0]) +
	( 2'sd 1) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_255;
assign conv_mac_255 = 
	( 3'sd 2) * $signed(input_fmap_1[7:0]) +
	( 2'sd 1) * $signed(input_fmap_2[7:0]) +
	( 2'sd 1) * $signed(input_fmap_3[7:0]) +
	( 2'sd 1) * $signed(input_fmap_6[7:0]) +
	( 3'sd 2) * $signed(input_fmap_7[7:0]) +
	( 2'sd 1) * $signed(input_fmap_8[7:0]) +
	( 2'sd 1) * $signed(input_fmap_10[7:0]) +
	( 2'sd 1) * $signed(input_fmap_11[7:0]) +
	( 2'sd 1) * $signed(input_fmap_12[7:0]) +
	( 2'sd 1) * $signed(input_fmap_16[7:0]) +
	( 2'sd 1) * $signed(input_fmap_17[7:0]) +
	( 3'sd 2) * $signed(input_fmap_18[7:0]) +
	( 3'sd 2) * $signed(input_fmap_20[7:0]) +
	( 2'sd 1) * $signed(input_fmap_22[7:0]) +
	( 2'sd 1) * $signed(input_fmap_23[7:0]) +
	( 2'sd 1) * $signed(input_fmap_24[7:0]) +
	( 2'sd 1) * $signed(input_fmap_25[7:0]) +
	( 2'sd 1) * $signed(input_fmap_26[7:0]) +
	( 2'sd 1) * $signed(input_fmap_27[7:0]) +
	( 2'sd 1) * $signed(input_fmap_28[7:0]) +
	( 2'sd 1) * $signed(input_fmap_29[7:0]) +
	( 2'sd 1) * $signed(input_fmap_31[7:0]) +
	( 2'sd 1) * $signed(input_fmap_32[7:0]) +
	( 2'sd 1) * $signed(input_fmap_35[7:0]) +
	( 3'sd 2) * $signed(input_fmap_37[7:0]) +
	( 2'sd 1) * $signed(input_fmap_38[7:0]) +
	( 2'sd 1) * $signed(input_fmap_39[7:0]) +
	( 2'sd 1) * $signed(input_fmap_40[7:0]) +
	( 3'sd 2) * $signed(input_fmap_41[7:0]) +
	( 2'sd 1) * $signed(input_fmap_42[7:0]) +
	( 3'sd 2) * $signed(input_fmap_43[7:0]) +
	( 2'sd 1) * $signed(input_fmap_44[7:0]) +
	( 3'sd 2) * $signed(input_fmap_45[7:0]) +
	( 2'sd 1) * $signed(input_fmap_48[7:0]) +
	( 2'sd 1) * $signed(input_fmap_50[7:0]) +
	( 2'sd 1) * $signed(input_fmap_51[7:0]) +
	( 2'sd 1) * $signed(input_fmap_54[7:0]) +
	( 2'sd 1) * $signed(input_fmap_56[7:0]) +
	( 2'sd 1) * $signed(input_fmap_57[7:0]) +
	( 2'sd 1) * $signed(input_fmap_58[7:0]) +
	( 2'sd 1) * $signed(input_fmap_59[7:0]) +
	( 2'sd 1) * $signed(input_fmap_62[7:0]) +
	( 2'sd 1) * $signed(input_fmap_63[7:0]) +
	( 2'sd 1) * $signed(input_fmap_64[7:0]) +
	( 3'sd 2) * $signed(input_fmap_66[7:0]) +
	( 2'sd 1) * $signed(input_fmap_67[7:0]) +
	( 2'sd 1) * $signed(input_fmap_69[7:0]) +
	( 2'sd 1) * $signed(input_fmap_70[7:0]) +
	( 2'sd 1) * $signed(input_fmap_72[7:0]) +
	( 2'sd 1) * $signed(input_fmap_73[7:0]) +
	( 2'sd 1) * $signed(input_fmap_74[7:0]) +
	( 3'sd 2) * $signed(input_fmap_75[7:0]) +
	( 2'sd 1) * $signed(input_fmap_76[7:0]) +
	( 2'sd 1) * $signed(input_fmap_77[7:0]) +
	( 3'sd 2) * $signed(input_fmap_78[7:0]) +
	( 2'sd 1) * $signed(input_fmap_79[7:0]) +
	( 2'sd 1) * $signed(input_fmap_80[7:0]) +
	( 2'sd 1) * $signed(input_fmap_81[7:0]) +
	( 3'sd 2) * $signed(input_fmap_82[7:0]) +
	( 2'sd 1) * $signed(input_fmap_83[7:0]) +
	( 2'sd 1) * $signed(input_fmap_84[7:0]) +
	( 2'sd 1) * $signed(input_fmap_85[7:0]) +
	( 2'sd 1) * $signed(input_fmap_86[7:0]) +
	( 2'sd 1) * $signed(input_fmap_87[7:0]) +
	( 3'sd 2) * $signed(input_fmap_89[7:0]) +
	( 3'sd 2) * $signed(input_fmap_91[7:0]) +
	( 3'sd 2) * $signed(input_fmap_94[7:0]) +
	( 3'sd 2) * $signed(input_fmap_95[7:0]) +
	( 2'sd 1) * $signed(input_fmap_96[7:0]) +
	( 2'sd 1) * $signed(input_fmap_97[7:0]) +
	( 2'sd 1) * $signed(input_fmap_98[7:0]) +
	( 3'sd 2) * $signed(input_fmap_99[7:0]) +
	( 2'sd 1) * $signed(input_fmap_100[7:0]) +
	( 2'sd 1) * $signed(input_fmap_101[7:0]) +
	( 2'sd 1) * $signed(input_fmap_102[7:0]) +
	( 2'sd 1) * $signed(input_fmap_103[7:0]) +
	( 3'sd 2) * $signed(input_fmap_104[7:0]) +
	( 2'sd 1) * $signed(input_fmap_105[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 2'sd 1) * $signed(input_fmap_111[7:0]) +
	( 3'sd 2) * $signed(input_fmap_112[7:0]) +
	( 3'sd 2) * $signed(input_fmap_114[7:0]) +
	( 3'sd 2) * $signed(input_fmap_116[7:0]) +
	( 2'sd 1) * $signed(input_fmap_117[7:0]) +
	( 3'sd 2) * $signed(input_fmap_118[7:0]) +
	( 2'sd 1) * $signed(input_fmap_119[7:0]) +
	( 2'sd 1) * $signed(input_fmap_120[7:0]) +
	( 2'sd 1) * $signed(input_fmap_121[7:0]) +
	( 2'sd 1) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 3'sd 2) * $signed(input_fmap_124[7:0]) +
	( 3'sd 2) * $signed(input_fmap_125[7:0]) +
	( 2'sd 1) * $signed(input_fmap_126[7:0]) +
	( 2'sd 1) * $signed(input_fmap_128[7:0]) +
	( 3'sd 2) * $signed(input_fmap_129[7:0]) +
	( 3'sd 2) * $signed(input_fmap_130[7:0]) +
	( 2'sd 1) * $signed(input_fmap_131[7:0]) +
	( 3'sd 2) * $signed(input_fmap_133[7:0]) +
	( 2'sd 1) * $signed(input_fmap_134[7:0]) +
	( 2'sd 1) * $signed(input_fmap_135[7:0]) +
	( 2'sd 1) * $signed(input_fmap_137[7:0]) +
	( 3'sd 2) * $signed(input_fmap_138[7:0]) +
	( 2'sd 1) * $signed(input_fmap_139[7:0]) +
	( 2'sd 1) * $signed(input_fmap_142[7:0]) +
	( 3'sd 2) * $signed(input_fmap_143[7:0]) +
	( 3'sd 2) * $signed(input_fmap_145[7:0]) +
	( 2'sd 1) * $signed(input_fmap_147[7:0]) +
	( 3'sd 2) * $signed(input_fmap_149[7:0]) +
	( 3'sd 2) * $signed(input_fmap_151[7:0]) +
	( 3'sd 2) * $signed(input_fmap_152[7:0]) +
	( 3'sd 2) * $signed(input_fmap_153[7:0]) +
	( 3'sd 2) * $signed(input_fmap_154[7:0]) +
	( 2'sd 1) * $signed(input_fmap_155[7:0]) +
	( 2'sd 1) * $signed(input_fmap_156[7:0]) +
	( 3'sd 2) * $signed(input_fmap_157[7:0]) +
	( 2'sd 1) * $signed(input_fmap_158[7:0]) +
	( 3'sd 2) * $signed(input_fmap_160[7:0]) +
	( 2'sd 1) * $signed(input_fmap_161[7:0]) +
	( 2'sd 1) * $signed(input_fmap_162[7:0]) +
	( 3'sd 2) * $signed(input_fmap_163[7:0]) +
	( 3'sd 2) * $signed(input_fmap_166[7:0]) +
	( 2'sd 1) * $signed(input_fmap_167[7:0]) +
	( 3'sd 2) * $signed(input_fmap_168[7:0]) +
	( 3'sd 2) * $signed(input_fmap_169[7:0]) +
	( 2'sd 1) * $signed(input_fmap_171[7:0]) +
	( 2'sd 1) * $signed(input_fmap_172[7:0]) +
	( 2'sd 1) * $signed(input_fmap_173[7:0]) +
	( 2'sd 1) * $signed(input_fmap_175[7:0]) +
	( 3'sd 2) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_178[7:0]) +
	( 2'sd 1) * $signed(input_fmap_179[7:0]) +
	( 2'sd 1) * $signed(input_fmap_180[7:0]) +
	( 2'sd 1) * $signed(input_fmap_181[7:0]) +
	( 2'sd 1) * $signed(input_fmap_182[7:0]) +
	( 2'sd 1) * $signed(input_fmap_183[7:0]) +
	( 3'sd 2) * $signed(input_fmap_185[7:0]) +
	( 2'sd 1) * $signed(input_fmap_186[7:0]) +
	( 2'sd 1) * $signed(input_fmap_188[7:0]) +
	( 3'sd 2) * $signed(input_fmap_189[7:0]) +
	( 2'sd 1) * $signed(input_fmap_192[7:0]) +
	( 3'sd 2) * $signed(input_fmap_193[7:0]) +
	( 2'sd 1) * $signed(input_fmap_195[7:0]) +
	( 2'sd 1) * $signed(input_fmap_196[7:0]) +
	( 2'sd 1) * $signed(input_fmap_197[7:0]) +
	( 3'sd 2) * $signed(input_fmap_199[7:0]) +
	( 2'sd 1) * $signed(input_fmap_200[7:0]) +
	( 2'sd 1) * $signed(input_fmap_203[7:0]) +
	( 2'sd 1) * $signed(input_fmap_204[7:0]) +
	( 2'sd 1) * $signed(input_fmap_205[7:0]) +
	( 3'sd 2) * $signed(input_fmap_206[7:0]) +
	( 2'sd 1) * $signed(input_fmap_207[7:0]) +
	( 3'sd 2) * $signed(input_fmap_208[7:0]) +
	( 2'sd 1) * $signed(input_fmap_210[7:0]) +
	( 3'sd 2) * $signed(input_fmap_211[7:0]) +
	( 2'sd 1) * $signed(input_fmap_212[7:0]) +
	( 3'sd 2) * $signed(input_fmap_214[7:0]) +
	( 2'sd 1) * $signed(input_fmap_217[7:0]) +
	( 2'sd 1) * $signed(input_fmap_219[7:0]) +
	( 2'sd 1) * $signed(input_fmap_221[7:0]) +
	( 3'sd 2) * $signed(input_fmap_222[7:0]) +
	( 2'sd 1) * $signed(input_fmap_223[7:0]) +
	( 2'sd 1) * $signed(input_fmap_225[7:0]) +
	( 2'sd 1) * $signed(input_fmap_230[7:0]) +
	( 2'sd 1) * $signed(input_fmap_231[7:0]) +
	( 2'sd 1) * $signed(input_fmap_232[7:0]) +
	( 2'sd 1) * $signed(input_fmap_234[7:0]) +
	( 3'sd 2) * $signed(input_fmap_235[7:0]) +
	( 2'sd 1) * $signed(input_fmap_237[7:0]) +
	( 2'sd 1) * $signed(input_fmap_238[7:0]) +
	( 2'sd 1) * $signed(input_fmap_239[7:0]) +
	( 2'sd 1) * $signed(input_fmap_241[7:0]) +
	( 2'sd 1) * $signed(input_fmap_242[7:0]) +
	( 2'sd 1) * $signed(input_fmap_243[7:0]) +
	( 3'sd 2) * $signed(input_fmap_244[7:0]) +
	( 2'sd 1) * $signed(input_fmap_245[7:0]) +
	( 2'sd 1) * $signed(input_fmap_246[7:0]) +
	( 2'sd 1) * $signed(input_fmap_247[7:0]) +
	( 3'sd 2) * $signed(input_fmap_249[7:0]) +
	( 3'sd 2) * $signed(input_fmap_252[7:0]) +
	( 3'sd 2) * $signed(input_fmap_253[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 3'd2;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 2'd1;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 2'd1;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 2'd1;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 2'd1;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 3'd2;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 2'd1;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 2'd1;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 2'd1;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 2'd1;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 3'd2;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 2'd1;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 3'd2;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 2'd1;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 2'd1;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 2'd1;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 2'd1;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 2'd1;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 2'd1;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 2'd1;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 2'd1;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 3'd2;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 3'd2;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 2'd1;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 2'd1;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 3'd2;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 2'd1;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 3'd2;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 2'd1;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 2'd1;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 2'd1;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 3'd2;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 2'd1;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 3'd2;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 2'd1;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 2'd1;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 3'd2;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 3'd2;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 2'd1;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 2'd1;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 3'd2;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 2'd1;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 3'd2;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 3'd2;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 2'd1;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 2'd1;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 2'd1;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 2'd1;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 2'd1;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 2'd1;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 2'd1;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 2'd1;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 2'd1;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 3'd2;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 3'd2;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 3'd2;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 2'd1;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 2'd1;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 2'd1;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 2'd1;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 2'd1;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 2'd1;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 2'd1;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 2'd1;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 2'd1;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 2'd1;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 2'd1;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 2'd1;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 3'd2;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 2'd1;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 2'd1;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 2'd1;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 2'd1;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 2'd1;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 2'd1;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 2'd1;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 2'd1;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 2'd1;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 3'd2;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 2'd1;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 3'd2;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 3'd2;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 2'd1;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 2'd1;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 2'd1;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 2'd1;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 3'd2;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 3'd2;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 2'd1;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 2'd1;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 2'd1;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 2'd1;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 2'd1;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 3'd2;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 2'd1;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 2'd1;
logic [31:0] bias_add_128;
assign bias_add_128 = conv_mac_128 + 2'd1;
logic [31:0] bias_add_129;
assign bias_add_129 = conv_mac_129 + 2'd1;
logic [31:0] bias_add_130;
assign bias_add_130 = conv_mac_130;
logic [31:0] bias_add_131;
assign bias_add_131 = conv_mac_131 + 2'd1;
logic [31:0] bias_add_132;
assign bias_add_132 = conv_mac_132 + 3'd2;
logic [31:0] bias_add_133;
assign bias_add_133 = conv_mac_133 + 2'd1;
logic [31:0] bias_add_134;
assign bias_add_134 = conv_mac_134 + 2'd1;
logic [31:0] bias_add_135;
assign bias_add_135 = conv_mac_135 + 3'd2;
logic [31:0] bias_add_136;
assign bias_add_136 = conv_mac_136 + 3'd2;
logic [31:0] bias_add_137;
assign bias_add_137 = conv_mac_137 + 3'd2;
logic [31:0] bias_add_138;
assign bias_add_138 = conv_mac_138 + 2'd1;
logic [31:0] bias_add_139;
assign bias_add_139 = conv_mac_139;
logic [31:0] bias_add_140;
assign bias_add_140 = conv_mac_140 + 2'd1;
logic [31:0] bias_add_141;
assign bias_add_141 = conv_mac_141;
logic [31:0] bias_add_142;
assign bias_add_142 = conv_mac_142;
logic [31:0] bias_add_143;
assign bias_add_143 = conv_mac_143 + 3'd2;
logic [31:0] bias_add_144;
assign bias_add_144 = conv_mac_144 + 2'd1;
logic [31:0] bias_add_145;
assign bias_add_145 = conv_mac_145 + 2'd1;
logic [31:0] bias_add_146;
assign bias_add_146 = conv_mac_146;
logic [31:0] bias_add_147;
assign bias_add_147 = conv_mac_147 + 3'd2;
logic [31:0] bias_add_148;
assign bias_add_148 = conv_mac_148 + 2'd1;
logic [31:0] bias_add_149;
assign bias_add_149 = conv_mac_149 + 3'd2;
logic [31:0] bias_add_150;
assign bias_add_150 = conv_mac_150;
logic [31:0] bias_add_151;
assign bias_add_151 = conv_mac_151 + 2'd1;
logic [31:0] bias_add_152;
assign bias_add_152 = conv_mac_152 + 2'd1;
logic [31:0] bias_add_153;
assign bias_add_153 = conv_mac_153 + 3'd2;
logic [31:0] bias_add_154;
assign bias_add_154 = conv_mac_154 + 2'd1;
logic [31:0] bias_add_155;
assign bias_add_155 = conv_mac_155 + 2'd1;
logic [31:0] bias_add_156;
assign bias_add_156 = conv_mac_156 + 3'd2;
logic [31:0] bias_add_157;
assign bias_add_157 = conv_mac_157;
logic [31:0] bias_add_158;
assign bias_add_158 = conv_mac_158 + 2'd1;
logic [31:0] bias_add_159;
assign bias_add_159 = conv_mac_159 + 2'd1;
logic [31:0] bias_add_160;
assign bias_add_160 = conv_mac_160 + 3'd2;
logic [31:0] bias_add_161;
assign bias_add_161 = conv_mac_161 + 2'd1;
logic [31:0] bias_add_162;
assign bias_add_162 = conv_mac_162 + 2'd1;
logic [31:0] bias_add_163;
assign bias_add_163 = conv_mac_163 + 3'd2;
logic [31:0] bias_add_164;
assign bias_add_164 = conv_mac_164 + 3'd2;
logic [31:0] bias_add_165;
assign bias_add_165 = conv_mac_165 + 3'd2;
logic [31:0] bias_add_166;
assign bias_add_166 = conv_mac_166;
logic [31:0] bias_add_167;
assign bias_add_167 = conv_mac_167 + 2'd1;
logic [31:0] bias_add_168;
assign bias_add_168 = conv_mac_168 + 2'd1;
logic [31:0] bias_add_169;
assign bias_add_169 = conv_mac_169 + 3'd2;
logic [31:0] bias_add_170;
assign bias_add_170 = conv_mac_170 + 2'd1;
logic [31:0] bias_add_171;
assign bias_add_171 = conv_mac_171 + 2'd1;
logic [31:0] bias_add_172;
assign bias_add_172 = conv_mac_172 + 3'd2;
logic [31:0] bias_add_173;
assign bias_add_173 = conv_mac_173 + 3'd2;
logic [31:0] bias_add_174;
assign bias_add_174 = conv_mac_174;
logic [31:0] bias_add_175;
assign bias_add_175 = conv_mac_175 + 3'd2;
logic [31:0] bias_add_176;
assign bias_add_176 = conv_mac_176 + 2'd1;
logic [31:0] bias_add_177;
assign bias_add_177 = conv_mac_177;
logic [31:0] bias_add_178;
assign bias_add_178 = conv_mac_178 + 2'd1;
logic [31:0] bias_add_179;
assign bias_add_179 = conv_mac_179 + 2'd1;
logic [31:0] bias_add_180;
assign bias_add_180 = conv_mac_180 + 2'd1;
logic [31:0] bias_add_181;
assign bias_add_181 = conv_mac_181 + 2'd1;
logic [31:0] bias_add_182;
assign bias_add_182 = conv_mac_182 + 2'd1;
logic [31:0] bias_add_183;
assign bias_add_183 = conv_mac_183 + 3'd2;
logic [31:0] bias_add_184;
assign bias_add_184 = conv_mac_184 + 2'd1;
logic [31:0] bias_add_185;
assign bias_add_185 = conv_mac_185 + 2'd1;
logic [31:0] bias_add_186;
assign bias_add_186 = conv_mac_186 + 2'd1;
logic [31:0] bias_add_187;
assign bias_add_187 = conv_mac_187 + 2'd1;
logic [31:0] bias_add_188;
assign bias_add_188 = conv_mac_188 + 3'd2;
logic [31:0] bias_add_189;
assign bias_add_189 = conv_mac_189;
logic [31:0] bias_add_190;
assign bias_add_190 = conv_mac_190;
logic [31:0] bias_add_191;
assign bias_add_191 = conv_mac_191;
logic [31:0] bias_add_192;
assign bias_add_192 = conv_mac_192 + 2'd1;
logic [31:0] bias_add_193;
assign bias_add_193 = conv_mac_193 + 2'd1;
logic [31:0] bias_add_194;
assign bias_add_194 = conv_mac_194 + 2'd1;
logic [31:0] bias_add_195;
assign bias_add_195 = conv_mac_195;
logic [31:0] bias_add_196;
assign bias_add_196 = conv_mac_196;
logic [31:0] bias_add_197;
assign bias_add_197 = conv_mac_197 + 3'd2;
logic [31:0] bias_add_198;
assign bias_add_198 = conv_mac_198 + 2'd1;
logic [31:0] bias_add_199;
assign bias_add_199 = conv_mac_199;
logic [31:0] bias_add_200;
assign bias_add_200 = conv_mac_200;
logic [31:0] bias_add_201;
assign bias_add_201 = conv_mac_201;
logic [31:0] bias_add_202;
assign bias_add_202 = conv_mac_202 + 3'd2;
logic [31:0] bias_add_203;
assign bias_add_203 = conv_mac_203;
logic [31:0] bias_add_204;
assign bias_add_204 = conv_mac_204 + 3'd2;
logic [31:0] bias_add_205;
assign bias_add_205 = conv_mac_205 + 2'd1;
logic [31:0] bias_add_206;
assign bias_add_206 = conv_mac_206 + 2'd1;
logic [31:0] bias_add_207;
assign bias_add_207 = conv_mac_207 + 2'd1;
logic [31:0] bias_add_208;
assign bias_add_208 = conv_mac_208 + 3'd2;
logic [31:0] bias_add_209;
assign bias_add_209 = conv_mac_209 + 2'd1;
logic [31:0] bias_add_210;
assign bias_add_210 = conv_mac_210 + 2'd1;
logic [31:0] bias_add_211;
assign bias_add_211 = conv_mac_211 + 3'd2;
logic [31:0] bias_add_212;
assign bias_add_212 = conv_mac_212;
logic [31:0] bias_add_213;
assign bias_add_213 = conv_mac_213 + 2'd1;
logic [31:0] bias_add_214;
assign bias_add_214 = conv_mac_214 + 2'd1;
logic [31:0] bias_add_215;
assign bias_add_215 = conv_mac_215 + 2'd1;
logic [31:0] bias_add_216;
assign bias_add_216 = conv_mac_216 + 3'd2;
logic [31:0] bias_add_217;
assign bias_add_217 = conv_mac_217;
logic [31:0] bias_add_218;
assign bias_add_218 = conv_mac_218 + 3'd2;
logic [31:0] bias_add_219;
assign bias_add_219 = conv_mac_219;
logic [31:0] bias_add_220;
assign bias_add_220 = conv_mac_220;
logic [31:0] bias_add_221;
assign bias_add_221 = conv_mac_221;
logic [31:0] bias_add_222;
assign bias_add_222 = conv_mac_222 + 2'd1;
logic [31:0] bias_add_223;
assign bias_add_223 = conv_mac_223;
logic [31:0] bias_add_224;
assign bias_add_224 = conv_mac_224 + 3'd2;
logic [31:0] bias_add_225;
assign bias_add_225 = conv_mac_225 + 3'd2;
logic [31:0] bias_add_226;
assign bias_add_226 = conv_mac_226 + 2'd1;
logic [31:0] bias_add_227;
assign bias_add_227 = conv_mac_227;
logic [31:0] bias_add_228;
assign bias_add_228 = conv_mac_228 + 2'd1;
logic [31:0] bias_add_229;
assign bias_add_229 = conv_mac_229;
logic [31:0] bias_add_230;
assign bias_add_230 = conv_mac_230 + 2'd1;
logic [31:0] bias_add_231;
assign bias_add_231 = conv_mac_231 + 3'd2;
logic [31:0] bias_add_232;
assign bias_add_232 = conv_mac_232 + 2'd1;
logic [31:0] bias_add_233;
assign bias_add_233 = conv_mac_233 + 3'd2;
logic [31:0] bias_add_234;
assign bias_add_234 = conv_mac_234;
logic [31:0] bias_add_235;
assign bias_add_235 = conv_mac_235 + 3'd2;
logic [31:0] bias_add_236;
assign bias_add_236 = conv_mac_236;
logic [31:0] bias_add_237;
assign bias_add_237 = conv_mac_237 + 3'd2;
logic [31:0] bias_add_238;
assign bias_add_238 = conv_mac_238;
logic [31:0] bias_add_239;
assign bias_add_239 = conv_mac_239 + 2'd1;
logic [31:0] bias_add_240;
assign bias_add_240 = conv_mac_240 + 3'd2;
logic [31:0] bias_add_241;
assign bias_add_241 = conv_mac_241;
logic [31:0] bias_add_242;
assign bias_add_242 = conv_mac_242 + 2'd1;
logic [31:0] bias_add_243;
assign bias_add_243 = conv_mac_243;
logic [31:0] bias_add_244;
assign bias_add_244 = conv_mac_244 + 3'd2;
logic [31:0] bias_add_245;
assign bias_add_245 = conv_mac_245 + 3'd2;
logic [31:0] bias_add_246;
assign bias_add_246 = conv_mac_246 + 2'd1;
logic [31:0] bias_add_247;
assign bias_add_247 = conv_mac_247 + 3'd2;
logic [31:0] bias_add_248;
assign bias_add_248 = conv_mac_248 + 2'd1;
logic [31:0] bias_add_249;
assign bias_add_249 = conv_mac_249 + 3'd2;
logic [31:0] bias_add_250;
assign bias_add_250 = conv_mac_250;
logic [31:0] bias_add_251;
assign bias_add_251 = conv_mac_251 + 3'd2;
logic [31:0] bias_add_252;
assign bias_add_252 = conv_mac_252 + 3'd2;
logic [31:0] bias_add_253;
assign bias_add_253 = conv_mac_253;
logic [31:0] bias_add_254;
assign bias_add_254 = conv_mac_254 + 2'd1;
logic [31:0] bias_add_255;
assign bias_add_255 = conv_mac_255;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[7:1]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[7:1]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[7:1]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[7:1]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[7:1]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[7:1]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[7:1]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[7:1]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[7:1]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[7:1]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[7:1]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[7:1]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[7:1]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[7:1]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[7:1]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[7:1]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[7:1]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[7:1]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[7:1]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[7:1]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[7:1]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[7:1]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[7:1]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[7:1]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[7:1]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[7:1]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[7:1]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[7:1]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[7:1]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[7:1]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[7:1]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[7:1]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[7:1]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[7:1]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[7:1]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[7:1]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[7:1]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[7:1]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[7:1]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[7:1]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[7:1]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[7:1]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[7:1]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[7:1]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[7:1]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[7:1]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[7:1]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[7:1]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[7:1]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[7:1]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[7:1]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[7:1]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[7:1]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[7:1]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[7:1]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[7:1]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[7:1]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[7:1]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[7:1]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[7:1]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[7:1]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[7:1]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[7:1]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[7:1]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[7:1]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[7:1]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[7:1]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[7:1]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[7:1]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[7:1]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[7:1]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[7:1]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[7:1]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[7:1]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[7:1]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[7:1]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[7:1]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[7:1]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[7:1]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[7:1]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[7:1]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[7:1]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[7:1]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[7:1]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[7:1]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[7:1]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[7:1]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[7:1]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[7:1]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[7:1]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[7:1]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[7:1]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[7:1]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[7:1]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[7:1]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[7:1]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[7:1]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[7:1]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[7:1]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[7:1]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[7:1]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[7:1]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[7:1]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[7:1]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[7:1]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[7:1]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[7:1]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[7:1]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[7:1]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[7:1]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[7:1]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[7:1]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[7:1]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[7:1]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[7:1]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[7:1]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[7:1]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[7:1]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[7:1]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[7:1]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[7:1]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[7:1]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[7:1]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[7:1]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[7:1]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[7:1]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[7:1]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[7:1]}} :'d6) : '0;
logic [7:0] relu_128;
assign relu_128[7:0] = (bias_add_128[31]==0) ? ((bias_add_128<3'd6) ? {{bias_add_128[31],bias_add_128[7:1]}} :'d6) : '0;
logic [7:0] relu_129;
assign relu_129[7:0] = (bias_add_129[31]==0) ? ((bias_add_129<3'd6) ? {{bias_add_129[31],bias_add_129[7:1]}} :'d6) : '0;
logic [7:0] relu_130;
assign relu_130[7:0] = (bias_add_130[31]==0) ? ((bias_add_130<3'd6) ? {{bias_add_130[31],bias_add_130[7:1]}} :'d6) : '0;
logic [7:0] relu_131;
assign relu_131[7:0] = (bias_add_131[31]==0) ? ((bias_add_131<3'd6) ? {{bias_add_131[31],bias_add_131[7:1]}} :'d6) : '0;
logic [7:0] relu_132;
assign relu_132[7:0] = (bias_add_132[31]==0) ? ((bias_add_132<3'd6) ? {{bias_add_132[31],bias_add_132[7:1]}} :'d6) : '0;
logic [7:0] relu_133;
assign relu_133[7:0] = (bias_add_133[31]==0) ? ((bias_add_133<3'd6) ? {{bias_add_133[31],bias_add_133[7:1]}} :'d6) : '0;
logic [7:0] relu_134;
assign relu_134[7:0] = (bias_add_134[31]==0) ? ((bias_add_134<3'd6) ? {{bias_add_134[31],bias_add_134[7:1]}} :'d6) : '0;
logic [7:0] relu_135;
assign relu_135[7:0] = (bias_add_135[31]==0) ? ((bias_add_135<3'd6) ? {{bias_add_135[31],bias_add_135[7:1]}} :'d6) : '0;
logic [7:0] relu_136;
assign relu_136[7:0] = (bias_add_136[31]==0) ? ((bias_add_136<3'd6) ? {{bias_add_136[31],bias_add_136[7:1]}} :'d6) : '0;
logic [7:0] relu_137;
assign relu_137[7:0] = (bias_add_137[31]==0) ? ((bias_add_137<3'd6) ? {{bias_add_137[31],bias_add_137[7:1]}} :'d6) : '0;
logic [7:0] relu_138;
assign relu_138[7:0] = (bias_add_138[31]==0) ? ((bias_add_138<3'd6) ? {{bias_add_138[31],bias_add_138[7:1]}} :'d6) : '0;
logic [7:0] relu_139;
assign relu_139[7:0] = (bias_add_139[31]==0) ? ((bias_add_139<3'd6) ? {{bias_add_139[31],bias_add_139[7:1]}} :'d6) : '0;
logic [7:0] relu_140;
assign relu_140[7:0] = (bias_add_140[31]==0) ? ((bias_add_140<3'd6) ? {{bias_add_140[31],bias_add_140[7:1]}} :'d6) : '0;
logic [7:0] relu_141;
assign relu_141[7:0] = (bias_add_141[31]==0) ? ((bias_add_141<3'd6) ? {{bias_add_141[31],bias_add_141[7:1]}} :'d6) : '0;
logic [7:0] relu_142;
assign relu_142[7:0] = (bias_add_142[31]==0) ? ((bias_add_142<3'd6) ? {{bias_add_142[31],bias_add_142[7:1]}} :'d6) : '0;
logic [7:0] relu_143;
assign relu_143[7:0] = (bias_add_143[31]==0) ? ((bias_add_143<3'd6) ? {{bias_add_143[31],bias_add_143[7:1]}} :'d6) : '0;
logic [7:0] relu_144;
assign relu_144[7:0] = (bias_add_144[31]==0) ? ((bias_add_144<3'd6) ? {{bias_add_144[31],bias_add_144[7:1]}} :'d6) : '0;
logic [7:0] relu_145;
assign relu_145[7:0] = (bias_add_145[31]==0) ? ((bias_add_145<3'd6) ? {{bias_add_145[31],bias_add_145[7:1]}} :'d6) : '0;
logic [7:0] relu_146;
assign relu_146[7:0] = (bias_add_146[31]==0) ? ((bias_add_146<3'd6) ? {{bias_add_146[31],bias_add_146[7:1]}} :'d6) : '0;
logic [7:0] relu_147;
assign relu_147[7:0] = (bias_add_147[31]==0) ? ((bias_add_147<3'd6) ? {{bias_add_147[31],bias_add_147[7:1]}} :'d6) : '0;
logic [7:0] relu_148;
assign relu_148[7:0] = (bias_add_148[31]==0) ? ((bias_add_148<3'd6) ? {{bias_add_148[31],bias_add_148[7:1]}} :'d6) : '0;
logic [7:0] relu_149;
assign relu_149[7:0] = (bias_add_149[31]==0) ? ((bias_add_149<3'd6) ? {{bias_add_149[31],bias_add_149[7:1]}} :'d6) : '0;
logic [7:0] relu_150;
assign relu_150[7:0] = (bias_add_150[31]==0) ? ((bias_add_150<3'd6) ? {{bias_add_150[31],bias_add_150[7:1]}} :'d6) : '0;
logic [7:0] relu_151;
assign relu_151[7:0] = (bias_add_151[31]==0) ? ((bias_add_151<3'd6) ? {{bias_add_151[31],bias_add_151[7:1]}} :'d6) : '0;
logic [7:0] relu_152;
assign relu_152[7:0] = (bias_add_152[31]==0) ? ((bias_add_152<3'd6) ? {{bias_add_152[31],bias_add_152[7:1]}} :'d6) : '0;
logic [7:0] relu_153;
assign relu_153[7:0] = (bias_add_153[31]==0) ? ((bias_add_153<3'd6) ? {{bias_add_153[31],bias_add_153[7:1]}} :'d6) : '0;
logic [7:0] relu_154;
assign relu_154[7:0] = (bias_add_154[31]==0) ? ((bias_add_154<3'd6) ? {{bias_add_154[31],bias_add_154[7:1]}} :'d6) : '0;
logic [7:0] relu_155;
assign relu_155[7:0] = (bias_add_155[31]==0) ? ((bias_add_155<3'd6) ? {{bias_add_155[31],bias_add_155[7:1]}} :'d6) : '0;
logic [7:0] relu_156;
assign relu_156[7:0] = (bias_add_156[31]==0) ? ((bias_add_156<3'd6) ? {{bias_add_156[31],bias_add_156[7:1]}} :'d6) : '0;
logic [7:0] relu_157;
assign relu_157[7:0] = (bias_add_157[31]==0) ? ((bias_add_157<3'd6) ? {{bias_add_157[31],bias_add_157[7:1]}} :'d6) : '0;
logic [7:0] relu_158;
assign relu_158[7:0] = (bias_add_158[31]==0) ? ((bias_add_158<3'd6) ? {{bias_add_158[31],bias_add_158[7:1]}} :'d6) : '0;
logic [7:0] relu_159;
assign relu_159[7:0] = (bias_add_159[31]==0) ? ((bias_add_159<3'd6) ? {{bias_add_159[31],bias_add_159[7:1]}} :'d6) : '0;
logic [7:0] relu_160;
assign relu_160[7:0] = (bias_add_160[31]==0) ? ((bias_add_160<3'd6) ? {{bias_add_160[31],bias_add_160[7:1]}} :'d6) : '0;
logic [7:0] relu_161;
assign relu_161[7:0] = (bias_add_161[31]==0) ? ((bias_add_161<3'd6) ? {{bias_add_161[31],bias_add_161[7:1]}} :'d6) : '0;
logic [7:0] relu_162;
assign relu_162[7:0] = (bias_add_162[31]==0) ? ((bias_add_162<3'd6) ? {{bias_add_162[31],bias_add_162[7:1]}} :'d6) : '0;
logic [7:0] relu_163;
assign relu_163[7:0] = (bias_add_163[31]==0) ? ((bias_add_163<3'd6) ? {{bias_add_163[31],bias_add_163[7:1]}} :'d6) : '0;
logic [7:0] relu_164;
assign relu_164[7:0] = (bias_add_164[31]==0) ? ((bias_add_164<3'd6) ? {{bias_add_164[31],bias_add_164[7:1]}} :'d6) : '0;
logic [7:0] relu_165;
assign relu_165[7:0] = (bias_add_165[31]==0) ? ((bias_add_165<3'd6) ? {{bias_add_165[31],bias_add_165[7:1]}} :'d6) : '0;
logic [7:0] relu_166;
assign relu_166[7:0] = (bias_add_166[31]==0) ? ((bias_add_166<3'd6) ? {{bias_add_166[31],bias_add_166[7:1]}} :'d6) : '0;
logic [7:0] relu_167;
assign relu_167[7:0] = (bias_add_167[31]==0) ? ((bias_add_167<3'd6) ? {{bias_add_167[31],bias_add_167[7:1]}} :'d6) : '0;
logic [7:0] relu_168;
assign relu_168[7:0] = (bias_add_168[31]==0) ? ((bias_add_168<3'd6) ? {{bias_add_168[31],bias_add_168[7:1]}} :'d6) : '0;
logic [7:0] relu_169;
assign relu_169[7:0] = (bias_add_169[31]==0) ? ((bias_add_169<3'd6) ? {{bias_add_169[31],bias_add_169[7:1]}} :'d6) : '0;
logic [7:0] relu_170;
assign relu_170[7:0] = (bias_add_170[31]==0) ? ((bias_add_170<3'd6) ? {{bias_add_170[31],bias_add_170[7:1]}} :'d6) : '0;
logic [7:0] relu_171;
assign relu_171[7:0] = (bias_add_171[31]==0) ? ((bias_add_171<3'd6) ? {{bias_add_171[31],bias_add_171[7:1]}} :'d6) : '0;
logic [7:0] relu_172;
assign relu_172[7:0] = (bias_add_172[31]==0) ? ((bias_add_172<3'd6) ? {{bias_add_172[31],bias_add_172[7:1]}} :'d6) : '0;
logic [7:0] relu_173;
assign relu_173[7:0] = (bias_add_173[31]==0) ? ((bias_add_173<3'd6) ? {{bias_add_173[31],bias_add_173[7:1]}} :'d6) : '0;
logic [7:0] relu_174;
assign relu_174[7:0] = (bias_add_174[31]==0) ? ((bias_add_174<3'd6) ? {{bias_add_174[31],bias_add_174[7:1]}} :'d6) : '0;
logic [7:0] relu_175;
assign relu_175[7:0] = (bias_add_175[31]==0) ? ((bias_add_175<3'd6) ? {{bias_add_175[31],bias_add_175[7:1]}} :'d6) : '0;
logic [7:0] relu_176;
assign relu_176[7:0] = (bias_add_176[31]==0) ? ((bias_add_176<3'd6) ? {{bias_add_176[31],bias_add_176[7:1]}} :'d6) : '0;
logic [7:0] relu_177;
assign relu_177[7:0] = (bias_add_177[31]==0) ? ((bias_add_177<3'd6) ? {{bias_add_177[31],bias_add_177[7:1]}} :'d6) : '0;
logic [7:0] relu_178;
assign relu_178[7:0] = (bias_add_178[31]==0) ? ((bias_add_178<3'd6) ? {{bias_add_178[31],bias_add_178[7:1]}} :'d6) : '0;
logic [7:0] relu_179;
assign relu_179[7:0] = (bias_add_179[31]==0) ? ((bias_add_179<3'd6) ? {{bias_add_179[31],bias_add_179[7:1]}} :'d6) : '0;
logic [7:0] relu_180;
assign relu_180[7:0] = (bias_add_180[31]==0) ? ((bias_add_180<3'd6) ? {{bias_add_180[31],bias_add_180[7:1]}} :'d6) : '0;
logic [7:0] relu_181;
assign relu_181[7:0] = (bias_add_181[31]==0) ? ((bias_add_181<3'd6) ? {{bias_add_181[31],bias_add_181[7:1]}} :'d6) : '0;
logic [7:0] relu_182;
assign relu_182[7:0] = (bias_add_182[31]==0) ? ((bias_add_182<3'd6) ? {{bias_add_182[31],bias_add_182[7:1]}} :'d6) : '0;
logic [7:0] relu_183;
assign relu_183[7:0] = (bias_add_183[31]==0) ? ((bias_add_183<3'd6) ? {{bias_add_183[31],bias_add_183[7:1]}} :'d6) : '0;
logic [7:0] relu_184;
assign relu_184[7:0] = (bias_add_184[31]==0) ? ((bias_add_184<3'd6) ? {{bias_add_184[31],bias_add_184[7:1]}} :'d6) : '0;
logic [7:0] relu_185;
assign relu_185[7:0] = (bias_add_185[31]==0) ? ((bias_add_185<3'd6) ? {{bias_add_185[31],bias_add_185[7:1]}} :'d6) : '0;
logic [7:0] relu_186;
assign relu_186[7:0] = (bias_add_186[31]==0) ? ((bias_add_186<3'd6) ? {{bias_add_186[31],bias_add_186[7:1]}} :'d6) : '0;
logic [7:0] relu_187;
assign relu_187[7:0] = (bias_add_187[31]==0) ? ((bias_add_187<3'd6) ? {{bias_add_187[31],bias_add_187[7:1]}} :'d6) : '0;
logic [7:0] relu_188;
assign relu_188[7:0] = (bias_add_188[31]==0) ? ((bias_add_188<3'd6) ? {{bias_add_188[31],bias_add_188[7:1]}} :'d6) : '0;
logic [7:0] relu_189;
assign relu_189[7:0] = (bias_add_189[31]==0) ? ((bias_add_189<3'd6) ? {{bias_add_189[31],bias_add_189[7:1]}} :'d6) : '0;
logic [7:0] relu_190;
assign relu_190[7:0] = (bias_add_190[31]==0) ? ((bias_add_190<3'd6) ? {{bias_add_190[31],bias_add_190[7:1]}} :'d6) : '0;
logic [7:0] relu_191;
assign relu_191[7:0] = (bias_add_191[31]==0) ? ((bias_add_191<3'd6) ? {{bias_add_191[31],bias_add_191[7:1]}} :'d6) : '0;
logic [7:0] relu_192;
assign relu_192[7:0] = (bias_add_192[31]==0) ? ((bias_add_192<3'd6) ? {{bias_add_192[31],bias_add_192[7:1]}} :'d6) : '0;
logic [7:0] relu_193;
assign relu_193[7:0] = (bias_add_193[31]==0) ? ((bias_add_193<3'd6) ? {{bias_add_193[31],bias_add_193[7:1]}} :'d6) : '0;
logic [7:0] relu_194;
assign relu_194[7:0] = (bias_add_194[31]==0) ? ((bias_add_194<3'd6) ? {{bias_add_194[31],bias_add_194[7:1]}} :'d6) : '0;
logic [7:0] relu_195;
assign relu_195[7:0] = (bias_add_195[31]==0) ? ((bias_add_195<3'd6) ? {{bias_add_195[31],bias_add_195[7:1]}} :'d6) : '0;
logic [7:0] relu_196;
assign relu_196[7:0] = (bias_add_196[31]==0) ? ((bias_add_196<3'd6) ? {{bias_add_196[31],bias_add_196[7:1]}} :'d6) : '0;
logic [7:0] relu_197;
assign relu_197[7:0] = (bias_add_197[31]==0) ? ((bias_add_197<3'd6) ? {{bias_add_197[31],bias_add_197[7:1]}} :'d6) : '0;
logic [7:0] relu_198;
assign relu_198[7:0] = (bias_add_198[31]==0) ? ((bias_add_198<3'd6) ? {{bias_add_198[31],bias_add_198[7:1]}} :'d6) : '0;
logic [7:0] relu_199;
assign relu_199[7:0] = (bias_add_199[31]==0) ? ((bias_add_199<3'd6) ? {{bias_add_199[31],bias_add_199[7:1]}} :'d6) : '0;
logic [7:0] relu_200;
assign relu_200[7:0] = (bias_add_200[31]==0) ? ((bias_add_200<3'd6) ? {{bias_add_200[31],bias_add_200[7:1]}} :'d6) : '0;
logic [7:0] relu_201;
assign relu_201[7:0] = (bias_add_201[31]==0) ? ((bias_add_201<3'd6) ? {{bias_add_201[31],bias_add_201[7:1]}} :'d6) : '0;
logic [7:0] relu_202;
assign relu_202[7:0] = (bias_add_202[31]==0) ? ((bias_add_202<3'd6) ? {{bias_add_202[31],bias_add_202[7:1]}} :'d6) : '0;
logic [7:0] relu_203;
assign relu_203[7:0] = (bias_add_203[31]==0) ? ((bias_add_203<3'd6) ? {{bias_add_203[31],bias_add_203[7:1]}} :'d6) : '0;
logic [7:0] relu_204;
assign relu_204[7:0] = (bias_add_204[31]==0) ? ((bias_add_204<3'd6) ? {{bias_add_204[31],bias_add_204[7:1]}} :'d6) : '0;
logic [7:0] relu_205;
assign relu_205[7:0] = (bias_add_205[31]==0) ? ((bias_add_205<3'd6) ? {{bias_add_205[31],bias_add_205[7:1]}} :'d6) : '0;
logic [7:0] relu_206;
assign relu_206[7:0] = (bias_add_206[31]==0) ? ((bias_add_206<3'd6) ? {{bias_add_206[31],bias_add_206[7:1]}} :'d6) : '0;
logic [7:0] relu_207;
assign relu_207[7:0] = (bias_add_207[31]==0) ? ((bias_add_207<3'd6) ? {{bias_add_207[31],bias_add_207[7:1]}} :'d6) : '0;
logic [7:0] relu_208;
assign relu_208[7:0] = (bias_add_208[31]==0) ? ((bias_add_208<3'd6) ? {{bias_add_208[31],bias_add_208[7:1]}} :'d6) : '0;
logic [7:0] relu_209;
assign relu_209[7:0] = (bias_add_209[31]==0) ? ((bias_add_209<3'd6) ? {{bias_add_209[31],bias_add_209[7:1]}} :'d6) : '0;
logic [7:0] relu_210;
assign relu_210[7:0] = (bias_add_210[31]==0) ? ((bias_add_210<3'd6) ? {{bias_add_210[31],bias_add_210[7:1]}} :'d6) : '0;
logic [7:0] relu_211;
assign relu_211[7:0] = (bias_add_211[31]==0) ? ((bias_add_211<3'd6) ? {{bias_add_211[31],bias_add_211[7:1]}} :'d6) : '0;
logic [7:0] relu_212;
assign relu_212[7:0] = (bias_add_212[31]==0) ? ((bias_add_212<3'd6) ? {{bias_add_212[31],bias_add_212[7:1]}} :'d6) : '0;
logic [7:0] relu_213;
assign relu_213[7:0] = (bias_add_213[31]==0) ? ((bias_add_213<3'd6) ? {{bias_add_213[31],bias_add_213[7:1]}} :'d6) : '0;
logic [7:0] relu_214;
assign relu_214[7:0] = (bias_add_214[31]==0) ? ((bias_add_214<3'd6) ? {{bias_add_214[31],bias_add_214[7:1]}} :'d6) : '0;
logic [7:0] relu_215;
assign relu_215[7:0] = (bias_add_215[31]==0) ? ((bias_add_215<3'd6) ? {{bias_add_215[31],bias_add_215[7:1]}} :'d6) : '0;
logic [7:0] relu_216;
assign relu_216[7:0] = (bias_add_216[31]==0) ? ((bias_add_216<3'd6) ? {{bias_add_216[31],bias_add_216[7:1]}} :'d6) : '0;
logic [7:0] relu_217;
assign relu_217[7:0] = (bias_add_217[31]==0) ? ((bias_add_217<3'd6) ? {{bias_add_217[31],bias_add_217[7:1]}} :'d6) : '0;
logic [7:0] relu_218;
assign relu_218[7:0] = (bias_add_218[31]==0) ? ((bias_add_218<3'd6) ? {{bias_add_218[31],bias_add_218[7:1]}} :'d6) : '0;
logic [7:0] relu_219;
assign relu_219[7:0] = (bias_add_219[31]==0) ? ((bias_add_219<3'd6) ? {{bias_add_219[31],bias_add_219[7:1]}} :'d6) : '0;
logic [7:0] relu_220;
assign relu_220[7:0] = (bias_add_220[31]==0) ? ((bias_add_220<3'd6) ? {{bias_add_220[31],bias_add_220[7:1]}} :'d6) : '0;
logic [7:0] relu_221;
assign relu_221[7:0] = (bias_add_221[31]==0) ? ((bias_add_221<3'd6) ? {{bias_add_221[31],bias_add_221[7:1]}} :'d6) : '0;
logic [7:0] relu_222;
assign relu_222[7:0] = (bias_add_222[31]==0) ? ((bias_add_222<3'd6) ? {{bias_add_222[31],bias_add_222[7:1]}} :'d6) : '0;
logic [7:0] relu_223;
assign relu_223[7:0] = (bias_add_223[31]==0) ? ((bias_add_223<3'd6) ? {{bias_add_223[31],bias_add_223[7:1]}} :'d6) : '0;
logic [7:0] relu_224;
assign relu_224[7:0] = (bias_add_224[31]==0) ? ((bias_add_224<3'd6) ? {{bias_add_224[31],bias_add_224[7:1]}} :'d6) : '0;
logic [7:0] relu_225;
assign relu_225[7:0] = (bias_add_225[31]==0) ? ((bias_add_225<3'd6) ? {{bias_add_225[31],bias_add_225[7:1]}} :'d6) : '0;
logic [7:0] relu_226;
assign relu_226[7:0] = (bias_add_226[31]==0) ? ((bias_add_226<3'd6) ? {{bias_add_226[31],bias_add_226[7:1]}} :'d6) : '0;
logic [7:0] relu_227;
assign relu_227[7:0] = (bias_add_227[31]==0) ? ((bias_add_227<3'd6) ? {{bias_add_227[31],bias_add_227[7:1]}} :'d6) : '0;
logic [7:0] relu_228;
assign relu_228[7:0] = (bias_add_228[31]==0) ? ((bias_add_228<3'd6) ? {{bias_add_228[31],bias_add_228[7:1]}} :'d6) : '0;
logic [7:0] relu_229;
assign relu_229[7:0] = (bias_add_229[31]==0) ? ((bias_add_229<3'd6) ? {{bias_add_229[31],bias_add_229[7:1]}} :'d6) : '0;
logic [7:0] relu_230;
assign relu_230[7:0] = (bias_add_230[31]==0) ? ((bias_add_230<3'd6) ? {{bias_add_230[31],bias_add_230[7:1]}} :'d6) : '0;
logic [7:0] relu_231;
assign relu_231[7:0] = (bias_add_231[31]==0) ? ((bias_add_231<3'd6) ? {{bias_add_231[31],bias_add_231[7:1]}} :'d6) : '0;
logic [7:0] relu_232;
assign relu_232[7:0] = (bias_add_232[31]==0) ? ((bias_add_232<3'd6) ? {{bias_add_232[31],bias_add_232[7:1]}} :'d6) : '0;
logic [7:0] relu_233;
assign relu_233[7:0] = (bias_add_233[31]==0) ? ((bias_add_233<3'd6) ? {{bias_add_233[31],bias_add_233[7:1]}} :'d6) : '0;
logic [7:0] relu_234;
assign relu_234[7:0] = (bias_add_234[31]==0) ? ((bias_add_234<3'd6) ? {{bias_add_234[31],bias_add_234[7:1]}} :'d6) : '0;
logic [7:0] relu_235;
assign relu_235[7:0] = (bias_add_235[31]==0) ? ((bias_add_235<3'd6) ? {{bias_add_235[31],bias_add_235[7:1]}} :'d6) : '0;
logic [7:0] relu_236;
assign relu_236[7:0] = (bias_add_236[31]==0) ? ((bias_add_236<3'd6) ? {{bias_add_236[31],bias_add_236[7:1]}} :'d6) : '0;
logic [7:0] relu_237;
assign relu_237[7:0] = (bias_add_237[31]==0) ? ((bias_add_237<3'd6) ? {{bias_add_237[31],bias_add_237[7:1]}} :'d6) : '0;
logic [7:0] relu_238;
assign relu_238[7:0] = (bias_add_238[31]==0) ? ((bias_add_238<3'd6) ? {{bias_add_238[31],bias_add_238[7:1]}} :'d6) : '0;
logic [7:0] relu_239;
assign relu_239[7:0] = (bias_add_239[31]==0) ? ((bias_add_239<3'd6) ? {{bias_add_239[31],bias_add_239[7:1]}} :'d6) : '0;
logic [7:0] relu_240;
assign relu_240[7:0] = (bias_add_240[31]==0) ? ((bias_add_240<3'd6) ? {{bias_add_240[31],bias_add_240[7:1]}} :'d6) : '0;
logic [7:0] relu_241;
assign relu_241[7:0] = (bias_add_241[31]==0) ? ((bias_add_241<3'd6) ? {{bias_add_241[31],bias_add_241[7:1]}} :'d6) : '0;
logic [7:0] relu_242;
assign relu_242[7:0] = (bias_add_242[31]==0) ? ((bias_add_242<3'd6) ? {{bias_add_242[31],bias_add_242[7:1]}} :'d6) : '0;
logic [7:0] relu_243;
assign relu_243[7:0] = (bias_add_243[31]==0) ? ((bias_add_243<3'd6) ? {{bias_add_243[31],bias_add_243[7:1]}} :'d6) : '0;
logic [7:0] relu_244;
assign relu_244[7:0] = (bias_add_244[31]==0) ? ((bias_add_244<3'd6) ? {{bias_add_244[31],bias_add_244[7:1]}} :'d6) : '0;
logic [7:0] relu_245;
assign relu_245[7:0] = (bias_add_245[31]==0) ? ((bias_add_245<3'd6) ? {{bias_add_245[31],bias_add_245[7:1]}} :'d6) : '0;
logic [7:0] relu_246;
assign relu_246[7:0] = (bias_add_246[31]==0) ? ((bias_add_246<3'd6) ? {{bias_add_246[31],bias_add_246[7:1]}} :'d6) : '0;
logic [7:0] relu_247;
assign relu_247[7:0] = (bias_add_247[31]==0) ? ((bias_add_247<3'd6) ? {{bias_add_247[31],bias_add_247[7:1]}} :'d6) : '0;
logic [7:0] relu_248;
assign relu_248[7:0] = (bias_add_248[31]==0) ? ((bias_add_248<3'd6) ? {{bias_add_248[31],bias_add_248[7:1]}} :'d6) : '0;
logic [7:0] relu_249;
assign relu_249[7:0] = (bias_add_249[31]==0) ? ((bias_add_249<3'd6) ? {{bias_add_249[31],bias_add_249[7:1]}} :'d6) : '0;
logic [7:0] relu_250;
assign relu_250[7:0] = (bias_add_250[31]==0) ? ((bias_add_250<3'd6) ? {{bias_add_250[31],bias_add_250[7:1]}} :'d6) : '0;
logic [7:0] relu_251;
assign relu_251[7:0] = (bias_add_251[31]==0) ? ((bias_add_251<3'd6) ? {{bias_add_251[31],bias_add_251[7:1]}} :'d6) : '0;
logic [7:0] relu_252;
assign relu_252[7:0] = (bias_add_252[31]==0) ? ((bias_add_252<3'd6) ? {{bias_add_252[31],bias_add_252[7:1]}} :'d6) : '0;
logic [7:0] relu_253;
assign relu_253[7:0] = (bias_add_253[31]==0) ? ((bias_add_253<3'd6) ? {{bias_add_253[31],bias_add_253[7:1]}} :'d6) : '0;
logic [7:0] relu_254;
assign relu_254[7:0] = (bias_add_254[31]==0) ? ((bias_add_254<3'd6) ? {{bias_add_254[31],bias_add_254[7:1]}} :'d6) : '0;
logic [7:0] relu_255;
assign relu_255[7:0] = (bias_add_255[31]==0) ? ((bias_add_255<3'd6) ? {{bias_add_255[31],bias_add_255[7:1]}} :'d6) : '0;

assign output_act = {
	relu_255,
	relu_254,
	relu_253,
	relu_252,
	relu_251,
	relu_250,
	relu_249,
	relu_248,
	relu_247,
	relu_246,
	relu_245,
	relu_244,
	relu_243,
	relu_242,
	relu_241,
	relu_240,
	relu_239,
	relu_238,
	relu_237,
	relu_236,
	relu_235,
	relu_234,
	relu_233,
	relu_232,
	relu_231,
	relu_230,
	relu_229,
	relu_228,
	relu_227,
	relu_226,
	relu_225,
	relu_224,
	relu_223,
	relu_222,
	relu_221,
	relu_220,
	relu_219,
	relu_218,
	relu_217,
	relu_216,
	relu_215,
	relu_214,
	relu_213,
	relu_212,
	relu_211,
	relu_210,
	relu_209,
	relu_208,
	relu_207,
	relu_206,
	relu_205,
	relu_204,
	relu_203,
	relu_202,
	relu_201,
	relu_200,
	relu_199,
	relu_198,
	relu_197,
	relu_196,
	relu_195,
	relu_194,
	relu_193,
	relu_192,
	relu_191,
	relu_190,
	relu_189,
	relu_188,
	relu_187,
	relu_186,
	relu_185,
	relu_184,
	relu_183,
	relu_182,
	relu_181,
	relu_180,
	relu_179,
	relu_178,
	relu_177,
	relu_176,
	relu_175,
	relu_174,
	relu_173,
	relu_172,
	relu_171,
	relu_170,
	relu_169,
	relu_168,
	relu_167,
	relu_166,
	relu_165,
	relu_164,
	relu_163,
	relu_162,
	relu_161,
	relu_160,
	relu_159,
	relu_158,
	relu_157,
	relu_156,
	relu_155,
	relu_154,
	relu_153,
	relu_152,
	relu_151,
	relu_150,
	relu_149,
	relu_148,
	relu_147,
	relu_146,
	relu_145,
	relu_144,
	relu_143,
	relu_142,
	relu_141,
	relu_140,
	relu_139,
	relu_138,
	relu_137,
	relu_136,
	relu_135,
	relu_134,
	relu_133,
	relu_132,
	relu_131,
	relu_130,
	relu_129,
	relu_128,
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
