module conv14_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [4096-1:0] input_act,
    output logic [4096-1:0] output_act,
    output logic ready
);

logic [4096-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [15:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[15:0];
logic [15:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[31:16];
logic [15:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[47:32];
logic [15:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[63:48];
logic [15:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[79:64];
logic [15:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[95:80];
logic [15:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[111:96];
logic [15:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[127:112];
logic [15:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[143:128];
logic [15:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[159:144];
logic [15:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[175:160];
logic [15:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[191:176];
logic [15:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[207:192];
logic [15:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[223:208];
logic [15:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[239:224];
logic [15:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[255:240];
logic [15:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[271:256];
logic [15:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[287:272];
logic [15:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[303:288];
logic [15:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[319:304];
logic [15:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[335:320];
logic [15:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[351:336];
logic [15:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[367:352];
logic [15:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[383:368];
logic [15:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[399:384];
logic [15:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[415:400];
logic [15:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[431:416];
logic [15:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[447:432];
logic [15:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[463:448];
logic [15:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[479:464];
logic [15:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[495:480];
logic [15:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[511:496];
logic [15:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[527:512];
logic [15:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[543:528];
logic [15:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[559:544];
logic [15:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[575:560];
logic [15:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[591:576];
logic [15:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[607:592];
logic [15:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[623:608];
logic [15:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[639:624];
logic [15:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[655:640];
logic [15:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[671:656];
logic [15:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[687:672];
logic [15:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[703:688];
logic [15:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[719:704];
logic [15:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[735:720];
logic [15:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[751:736];
logic [15:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[767:752];
logic [15:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[783:768];
logic [15:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[799:784];
logic [15:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[815:800];
logic [15:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[831:816];
logic [15:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[847:832];
logic [15:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[863:848];
logic [15:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[879:864];
logic [15:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[895:880];
logic [15:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[911:896];
logic [15:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[927:912];
logic [15:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[943:928];
logic [15:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[959:944];
logic [15:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[975:960];
logic [15:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[991:976];
logic [15:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[1007:992];
logic [15:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[1023:1008];
logic [15:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[1039:1024];
logic [15:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[1055:1040];
logic [15:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[1071:1056];
logic [15:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[1087:1072];
logic [15:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[1103:1088];
logic [15:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[1119:1104];
logic [15:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[1135:1120];
logic [15:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[1151:1136];
logic [15:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[1167:1152];
logic [15:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[1183:1168];
logic [15:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[1199:1184];
logic [15:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[1215:1200];
logic [15:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[1231:1216];
logic [15:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[1247:1232];
logic [15:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[1263:1248];
logic [15:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[1279:1264];
logic [15:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[1295:1280];
logic [15:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[1311:1296];
logic [15:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[1327:1312];
logic [15:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[1343:1328];
logic [15:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[1359:1344];
logic [15:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[1375:1360];
logic [15:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[1391:1376];
logic [15:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[1407:1392];
logic [15:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[1423:1408];
logic [15:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[1439:1424];
logic [15:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[1455:1440];
logic [15:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[1471:1456];
logic [15:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[1487:1472];
logic [15:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[1503:1488];
logic [15:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[1519:1504];
logic [15:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[1535:1520];
logic [15:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[1551:1536];
logic [15:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[1567:1552];
logic [15:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[1583:1568];
logic [15:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[1599:1584];
logic [15:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[1615:1600];
logic [15:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[1631:1616];
logic [15:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[1647:1632];
logic [15:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[1663:1648];
logic [15:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[1679:1664];
logic [15:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[1695:1680];
logic [15:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[1711:1696];
logic [15:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[1727:1712];
logic [15:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[1743:1728];
logic [15:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[1759:1744];
logic [15:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[1775:1760];
logic [15:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[1791:1776];
logic [15:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[1807:1792];
logic [15:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[1823:1808];
logic [15:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[1839:1824];
logic [15:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[1855:1840];
logic [15:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[1871:1856];
logic [15:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[1887:1872];
logic [15:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[1903:1888];
logic [15:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[1919:1904];
logic [15:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[1935:1920];
logic [15:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[1951:1936];
logic [15:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[1967:1952];
logic [15:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[1983:1968];
logic [15:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[1999:1984];
logic [15:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[2015:2000];
logic [15:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[2031:2016];
logic [15:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[2047:2032];
logic [15:0] input_fmap_128;
assign input_fmap_128 = input_act_ff[2063:2048];
logic [15:0] input_fmap_129;
assign input_fmap_129 = input_act_ff[2079:2064];
logic [15:0] input_fmap_130;
assign input_fmap_130 = input_act_ff[2095:2080];
logic [15:0] input_fmap_131;
assign input_fmap_131 = input_act_ff[2111:2096];
logic [15:0] input_fmap_132;
assign input_fmap_132 = input_act_ff[2127:2112];
logic [15:0] input_fmap_133;
assign input_fmap_133 = input_act_ff[2143:2128];
logic [15:0] input_fmap_134;
assign input_fmap_134 = input_act_ff[2159:2144];
logic [15:0] input_fmap_135;
assign input_fmap_135 = input_act_ff[2175:2160];
logic [15:0] input_fmap_136;
assign input_fmap_136 = input_act_ff[2191:2176];
logic [15:0] input_fmap_137;
assign input_fmap_137 = input_act_ff[2207:2192];
logic [15:0] input_fmap_138;
assign input_fmap_138 = input_act_ff[2223:2208];
logic [15:0] input_fmap_139;
assign input_fmap_139 = input_act_ff[2239:2224];
logic [15:0] input_fmap_140;
assign input_fmap_140 = input_act_ff[2255:2240];
logic [15:0] input_fmap_141;
assign input_fmap_141 = input_act_ff[2271:2256];
logic [15:0] input_fmap_142;
assign input_fmap_142 = input_act_ff[2287:2272];
logic [15:0] input_fmap_143;
assign input_fmap_143 = input_act_ff[2303:2288];
logic [15:0] input_fmap_144;
assign input_fmap_144 = input_act_ff[2319:2304];
logic [15:0] input_fmap_145;
assign input_fmap_145 = input_act_ff[2335:2320];
logic [15:0] input_fmap_146;
assign input_fmap_146 = input_act_ff[2351:2336];
logic [15:0] input_fmap_147;
assign input_fmap_147 = input_act_ff[2367:2352];
logic [15:0] input_fmap_148;
assign input_fmap_148 = input_act_ff[2383:2368];
logic [15:0] input_fmap_149;
assign input_fmap_149 = input_act_ff[2399:2384];
logic [15:0] input_fmap_150;
assign input_fmap_150 = input_act_ff[2415:2400];
logic [15:0] input_fmap_151;
assign input_fmap_151 = input_act_ff[2431:2416];
logic [15:0] input_fmap_152;
assign input_fmap_152 = input_act_ff[2447:2432];
logic [15:0] input_fmap_153;
assign input_fmap_153 = input_act_ff[2463:2448];
logic [15:0] input_fmap_154;
assign input_fmap_154 = input_act_ff[2479:2464];
logic [15:0] input_fmap_155;
assign input_fmap_155 = input_act_ff[2495:2480];
logic [15:0] input_fmap_156;
assign input_fmap_156 = input_act_ff[2511:2496];
logic [15:0] input_fmap_157;
assign input_fmap_157 = input_act_ff[2527:2512];
logic [15:0] input_fmap_158;
assign input_fmap_158 = input_act_ff[2543:2528];
logic [15:0] input_fmap_159;
assign input_fmap_159 = input_act_ff[2559:2544];
logic [15:0] input_fmap_160;
assign input_fmap_160 = input_act_ff[2575:2560];
logic [15:0] input_fmap_161;
assign input_fmap_161 = input_act_ff[2591:2576];
logic [15:0] input_fmap_162;
assign input_fmap_162 = input_act_ff[2607:2592];
logic [15:0] input_fmap_163;
assign input_fmap_163 = input_act_ff[2623:2608];
logic [15:0] input_fmap_164;
assign input_fmap_164 = input_act_ff[2639:2624];
logic [15:0] input_fmap_165;
assign input_fmap_165 = input_act_ff[2655:2640];
logic [15:0] input_fmap_166;
assign input_fmap_166 = input_act_ff[2671:2656];
logic [15:0] input_fmap_167;
assign input_fmap_167 = input_act_ff[2687:2672];
logic [15:0] input_fmap_168;
assign input_fmap_168 = input_act_ff[2703:2688];
logic [15:0] input_fmap_169;
assign input_fmap_169 = input_act_ff[2719:2704];
logic [15:0] input_fmap_170;
assign input_fmap_170 = input_act_ff[2735:2720];
logic [15:0] input_fmap_171;
assign input_fmap_171 = input_act_ff[2751:2736];
logic [15:0] input_fmap_172;
assign input_fmap_172 = input_act_ff[2767:2752];
logic [15:0] input_fmap_173;
assign input_fmap_173 = input_act_ff[2783:2768];
logic [15:0] input_fmap_174;
assign input_fmap_174 = input_act_ff[2799:2784];
logic [15:0] input_fmap_175;
assign input_fmap_175 = input_act_ff[2815:2800];
logic [15:0] input_fmap_176;
assign input_fmap_176 = input_act_ff[2831:2816];
logic [15:0] input_fmap_177;
assign input_fmap_177 = input_act_ff[2847:2832];
logic [15:0] input_fmap_178;
assign input_fmap_178 = input_act_ff[2863:2848];
logic [15:0] input_fmap_179;
assign input_fmap_179 = input_act_ff[2879:2864];
logic [15:0] input_fmap_180;
assign input_fmap_180 = input_act_ff[2895:2880];
logic [15:0] input_fmap_181;
assign input_fmap_181 = input_act_ff[2911:2896];
logic [15:0] input_fmap_182;
assign input_fmap_182 = input_act_ff[2927:2912];
logic [15:0] input_fmap_183;
assign input_fmap_183 = input_act_ff[2943:2928];
logic [15:0] input_fmap_184;
assign input_fmap_184 = input_act_ff[2959:2944];
logic [15:0] input_fmap_185;
assign input_fmap_185 = input_act_ff[2975:2960];
logic [15:0] input_fmap_186;
assign input_fmap_186 = input_act_ff[2991:2976];
logic [15:0] input_fmap_187;
assign input_fmap_187 = input_act_ff[3007:2992];
logic [15:0] input_fmap_188;
assign input_fmap_188 = input_act_ff[3023:3008];
logic [15:0] input_fmap_189;
assign input_fmap_189 = input_act_ff[3039:3024];
logic [15:0] input_fmap_190;
assign input_fmap_190 = input_act_ff[3055:3040];
logic [15:0] input_fmap_191;
assign input_fmap_191 = input_act_ff[3071:3056];
logic [15:0] input_fmap_192;
assign input_fmap_192 = input_act_ff[3087:3072];
logic [15:0] input_fmap_193;
assign input_fmap_193 = input_act_ff[3103:3088];
logic [15:0] input_fmap_194;
assign input_fmap_194 = input_act_ff[3119:3104];
logic [15:0] input_fmap_195;
assign input_fmap_195 = input_act_ff[3135:3120];
logic [15:0] input_fmap_196;
assign input_fmap_196 = input_act_ff[3151:3136];
logic [15:0] input_fmap_197;
assign input_fmap_197 = input_act_ff[3167:3152];
logic [15:0] input_fmap_198;
assign input_fmap_198 = input_act_ff[3183:3168];
logic [15:0] input_fmap_199;
assign input_fmap_199 = input_act_ff[3199:3184];
logic [15:0] input_fmap_200;
assign input_fmap_200 = input_act_ff[3215:3200];
logic [15:0] input_fmap_201;
assign input_fmap_201 = input_act_ff[3231:3216];
logic [15:0] input_fmap_202;
assign input_fmap_202 = input_act_ff[3247:3232];
logic [15:0] input_fmap_203;
assign input_fmap_203 = input_act_ff[3263:3248];
logic [15:0] input_fmap_204;
assign input_fmap_204 = input_act_ff[3279:3264];
logic [15:0] input_fmap_205;
assign input_fmap_205 = input_act_ff[3295:3280];
logic [15:0] input_fmap_206;
assign input_fmap_206 = input_act_ff[3311:3296];
logic [15:0] input_fmap_207;
assign input_fmap_207 = input_act_ff[3327:3312];
logic [15:0] input_fmap_208;
assign input_fmap_208 = input_act_ff[3343:3328];
logic [15:0] input_fmap_209;
assign input_fmap_209 = input_act_ff[3359:3344];
logic [15:0] input_fmap_210;
assign input_fmap_210 = input_act_ff[3375:3360];
logic [15:0] input_fmap_211;
assign input_fmap_211 = input_act_ff[3391:3376];
logic [15:0] input_fmap_212;
assign input_fmap_212 = input_act_ff[3407:3392];
logic [15:0] input_fmap_213;
assign input_fmap_213 = input_act_ff[3423:3408];
logic [15:0] input_fmap_214;
assign input_fmap_214 = input_act_ff[3439:3424];
logic [15:0] input_fmap_215;
assign input_fmap_215 = input_act_ff[3455:3440];
logic [15:0] input_fmap_216;
assign input_fmap_216 = input_act_ff[3471:3456];
logic [15:0] input_fmap_217;
assign input_fmap_217 = input_act_ff[3487:3472];
logic [15:0] input_fmap_218;
assign input_fmap_218 = input_act_ff[3503:3488];
logic [15:0] input_fmap_219;
assign input_fmap_219 = input_act_ff[3519:3504];
logic [15:0] input_fmap_220;
assign input_fmap_220 = input_act_ff[3535:3520];
logic [15:0] input_fmap_221;
assign input_fmap_221 = input_act_ff[3551:3536];
logic [15:0] input_fmap_222;
assign input_fmap_222 = input_act_ff[3567:3552];
logic [15:0] input_fmap_223;
assign input_fmap_223 = input_act_ff[3583:3568];
logic [15:0] input_fmap_224;
assign input_fmap_224 = input_act_ff[3599:3584];
logic [15:0] input_fmap_225;
assign input_fmap_225 = input_act_ff[3615:3600];
logic [15:0] input_fmap_226;
assign input_fmap_226 = input_act_ff[3631:3616];
logic [15:0] input_fmap_227;
assign input_fmap_227 = input_act_ff[3647:3632];
logic [15:0] input_fmap_228;
assign input_fmap_228 = input_act_ff[3663:3648];
logic [15:0] input_fmap_229;
assign input_fmap_229 = input_act_ff[3679:3664];
logic [15:0] input_fmap_230;
assign input_fmap_230 = input_act_ff[3695:3680];
logic [15:0] input_fmap_231;
assign input_fmap_231 = input_act_ff[3711:3696];
logic [15:0] input_fmap_232;
assign input_fmap_232 = input_act_ff[3727:3712];
logic [15:0] input_fmap_233;
assign input_fmap_233 = input_act_ff[3743:3728];
logic [15:0] input_fmap_234;
assign input_fmap_234 = input_act_ff[3759:3744];
logic [15:0] input_fmap_235;
assign input_fmap_235 = input_act_ff[3775:3760];
logic [15:0] input_fmap_236;
assign input_fmap_236 = input_act_ff[3791:3776];
logic [15:0] input_fmap_237;
assign input_fmap_237 = input_act_ff[3807:3792];
logic [15:0] input_fmap_238;
assign input_fmap_238 = input_act_ff[3823:3808];
logic [15:0] input_fmap_239;
assign input_fmap_239 = input_act_ff[3839:3824];
logic [15:0] input_fmap_240;
assign input_fmap_240 = input_act_ff[3855:3840];
logic [15:0] input_fmap_241;
assign input_fmap_241 = input_act_ff[3871:3856];
logic [15:0] input_fmap_242;
assign input_fmap_242 = input_act_ff[3887:3872];
logic [15:0] input_fmap_243;
assign input_fmap_243 = input_act_ff[3903:3888];
logic [15:0] input_fmap_244;
assign input_fmap_244 = input_act_ff[3919:3904];
logic [15:0] input_fmap_245;
assign input_fmap_245 = input_act_ff[3935:3920];
logic [15:0] input_fmap_246;
assign input_fmap_246 = input_act_ff[3951:3936];
logic [15:0] input_fmap_247;
assign input_fmap_247 = input_act_ff[3967:3952];
logic [15:0] input_fmap_248;
assign input_fmap_248 = input_act_ff[3983:3968];
logic [15:0] input_fmap_249;
assign input_fmap_249 = input_act_ff[3999:3984];
logic [15:0] input_fmap_250;
assign input_fmap_250 = input_act_ff[4015:4000];
logic [15:0] input_fmap_251;
assign input_fmap_251 = input_act_ff[4031:4016];
logic [15:0] input_fmap_252;
assign input_fmap_252 = input_act_ff[4047:4032];
logic [15:0] input_fmap_253;
assign input_fmap_253 = input_act_ff[4063:4048];
logic [15:0] input_fmap_254;
assign input_fmap_254 = input_act_ff[4079:4064];
logic [15:0] input_fmap_255;
assign input_fmap_255 = input_act_ff[4095:4080];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 5'sd 8) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 5'sd 8) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_128;
assign conv_mac_128 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_129;
assign conv_mac_129 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_130;
assign conv_mac_130 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_131;
assign conv_mac_131 = 
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_132;
assign conv_mac_132 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_133;
assign conv_mac_133 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_134;
assign conv_mac_134 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_135;
assign conv_mac_135 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_136;
assign conv_mac_136 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_137;
assign conv_mac_137 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_138;
assign conv_mac_138 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_139;
assign conv_mac_139 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_140;
assign conv_mac_140 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_141;
assign conv_mac_141 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_142;
assign conv_mac_142 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_143;
assign conv_mac_143 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_144;
assign conv_mac_144 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_145;
assign conv_mac_145 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_146;
assign conv_mac_146 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_147;
assign conv_mac_147 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_148;
assign conv_mac_148 = 
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_149;
assign conv_mac_149 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_150;
assign conv_mac_150 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_151;
assign conv_mac_151 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_152;
assign conv_mac_152 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_153;
assign conv_mac_153 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_154;
assign conv_mac_154 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_155;
assign conv_mac_155 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_156;
assign conv_mac_156 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 5'sd 8) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_157;
assign conv_mac_157 = 
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_158;
assign conv_mac_158 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_159;
assign conv_mac_159 = 
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_160;
assign conv_mac_160 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_161;
assign conv_mac_161 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_162;
assign conv_mac_162 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_163;
assign conv_mac_163 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_164;
assign conv_mac_164 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_165;
assign conv_mac_165 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_166;
assign conv_mac_166 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_167;
assign conv_mac_167 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_168;
assign conv_mac_168 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_169;
assign conv_mac_169 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_170;
assign conv_mac_170 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_171;
assign conv_mac_171 = 
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_172;
assign conv_mac_172 = 
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_173;
assign conv_mac_173 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 5'sd 8) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_174;
assign conv_mac_174 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_175;
assign conv_mac_175 = 
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_176;
assign conv_mac_176 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_177;
assign conv_mac_177 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_178;
assign conv_mac_178 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_179;
assign conv_mac_179 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_180;
assign conv_mac_180 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_181;
assign conv_mac_181 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_182;
assign conv_mac_182 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_183;
assign conv_mac_183 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_184;
assign conv_mac_184 = 
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_185;
assign conv_mac_185 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_186;
assign conv_mac_186 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_187;
assign conv_mac_187 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_188;
assign conv_mac_188 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_189;
assign conv_mac_189 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_190;
assign conv_mac_190 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_191;
assign conv_mac_191 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_192;
assign conv_mac_192 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 5'sd 8) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_193;
assign conv_mac_193 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_194;
assign conv_mac_194 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_195;
assign conv_mac_195 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_196;
assign conv_mac_196 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_197;
assign conv_mac_197 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_198;
assign conv_mac_198 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_199;
assign conv_mac_199 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 5'sd 8) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_200;
assign conv_mac_200 = 
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 5'sd 8) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 5'sd 8) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_201;
assign conv_mac_201 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 5'sd 8) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_202;
assign conv_mac_202 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 4) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_203;
assign conv_mac_203 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 5'sd 8) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_204;
assign conv_mac_204 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_205;
assign conv_mac_205 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_206;
assign conv_mac_206 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 5'sd 8) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_207;
assign conv_mac_207 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_208;
assign conv_mac_208 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_209;
assign conv_mac_209 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_210;
assign conv_mac_210 = 
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_211;
assign conv_mac_211 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_212;
assign conv_mac_212 = 
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 3'sd 3) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 5) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 5'sd 8) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_213;
assign conv_mac_213 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_214;
assign conv_mac_214 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 5'sd 8) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_215;
assign conv_mac_215 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 2'sd 1) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_216;
assign conv_mac_216 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 3) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_217;
assign conv_mac_217 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 4'sd 4) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 5'sd 8) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_218;
assign conv_mac_218 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_219;
assign conv_mac_219 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 5'sd 8) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 3'sd 2) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 5'sd 8) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 3'sd 2) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_220;
assign conv_mac_220 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 5'sd 8) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 5'sd 8) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 4) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 5'sd 8) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 4) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 5'sd 8) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_221;
assign conv_mac_221 = 
	( 3'sd 3) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 5'sd 8) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 5) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 5'sd 8) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_222;
assign conv_mac_222 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 5'sd 8) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 5'sd 8) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 5'sd 8) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 3) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_223;
assign conv_mac_223 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 5'sd 8) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 5'sd 8) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 5'sd 8) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 3'sd 3) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 5'sd 8) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_224;
assign conv_mac_224 = 
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 5) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 2) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 6) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 4) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 3'sd 3) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_225;
assign conv_mac_225 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 5'sd 8) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 5'sd 8) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 6) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 3'sd 3) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 5'sd 8) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 6) * $signed(input_fmap_166[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_226;
assign conv_mac_226 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 5'sd 8) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 5'sd 8) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 5'sd 8) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 2) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 4'sd 7) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 5'sd 8) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_227;
assign conv_mac_227 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 5'sd 8) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 5'sd 8) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 2'sd 1) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 5'sd 8) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 4) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 5'sd 8) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 5'sd 8) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 5) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_228;
assign conv_mac_228 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 2'sd 1) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 5) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 2'sd 1) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 5'sd 8) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 6) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 5'sd 8) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 3'sd 2) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 7) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 2) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_229;
assign conv_mac_229 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 5'sd 8) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 4'sd 7) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 5'sd 8) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 5) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 3'sd 2) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 2'sd 1) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 5'sd 8) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_230;
assign conv_mac_230 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 5'sd 8) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 5'sd 8) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 5'sd 8) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 2'sd 1) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 3'sd 3) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 3'sd 3) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 5'sd 8) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 2'sd 1) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 4) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 2'sd 1) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 2'sd 1) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 2'sd 1) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 2'sd 1) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_231;
assign conv_mac_231 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 4'sd 4) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 5'sd 8) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 6) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 3'sd 2) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 4'sd 5) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 4) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_232;
assign conv_mac_232 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 3'sd 2) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 2) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 3'sd 3) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 4) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 4'sd 6) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 5'sd 8) * $signed(input_fmap_122[15:0]) +
	( 5'sd 8) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 2'sd 1) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 4'sd 7) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 5'sd 8) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 7) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_233;
assign conv_mac_233 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 6) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 4) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 4'sd 5) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 7) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 7) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 3'sd 3) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 2'sd 1) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 5'sd 8) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_234;
assign conv_mac_234 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 2'sd 1) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 5'sd 8) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 3'sd 2) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_99[15:0]) +
	( 4'sd 5) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 5'sd 8) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 5'sd 8) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 3'sd 3) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 4'sd 6) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 5'sd 8) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 4'sd 6) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 4'sd 5) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 4'sd 5) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 4'sd 4) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 2) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 5'sd 8) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_235;
assign conv_mac_235 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 6) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 5'sd 8) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 5'sd 8) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 3'sd 2) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 5'sd 8) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 2) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 5'sd 8) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 2'sd 1) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 3'sd 3) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 6) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 4'sd 6) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 4) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 4) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 4) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 2'sd 1) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 6) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_236;
assign conv_mac_236 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 5'sd 8) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 2'sd 1) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 4'sd 5) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 5'sd 8) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 5'sd 8) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 2'sd 1) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 3'sd 3) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 4) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 3'sd 2) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 4'sd 6) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 5'sd 8) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 3'sd 3) * $signed(input_fmap_243[15:0]) +
	( 3'sd 2) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 5'sd 8) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 2'sd 1) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_237;
assign conv_mac_237 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 4) * $signed(input_fmap_6[15:0]) +
	( 5'sd 8) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 4'sd 6) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 2'sd 1) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 3'sd 2) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 2'sd 1) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 3) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 4'sd 4) * $signed(input_fmap_75[15:0]) +
	( 4'sd 5) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 5'sd 8) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 3'sd 3) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 3'sd 2) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 5) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_132[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 3'sd 2) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_151[15:0]) +
	( 4'sd 7) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 3'sd 2) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 5'sd 8) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 2'sd 1) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 5'sd 8) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 7) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 6) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_238;
assign conv_mac_238 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 5) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 4'sd 7) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 6) * $signed(input_fmap_27[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 7) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 5) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 4) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 5'sd 8) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 4'sd 5) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 5'sd 8) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 3) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 5) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 5) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 6) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 6) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 5) * $signed(input_fmap_215[15:0]) +
	( 4'sd 7) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 5'sd 8) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 6) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 5'sd 8) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_239;
assign conv_mac_239 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 4) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 7) * $signed(input_fmap_4[15:0]) +
	( 2'sd 1) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 2'sd 1) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 4'sd 7) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 4) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 4'sd 7) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 2'sd 1) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 4) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 3) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_65[15:0]) +
	( 4'sd 5) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 6) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 5) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_112[15:0]) +
	( 4'sd 7) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 5'sd 8) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 3) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 5'sd 8) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 5'sd 8) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 4'sd 4) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 6) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 4) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 2'sd 1) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 6) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 3'sd 3) * $signed(input_fmap_222[15:0]) +
	( 5'sd 8) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 4'sd 4) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 3'sd 2) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_240;
assign conv_mac_240 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 4'sd 6) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 2) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 4) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 5) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 5'sd 8) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 4'sd 7) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 5'sd 8) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 2'sd 1) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 4'sd 5) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 5'sd 8) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 6) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 7) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 2'sd 1) * $signed(input_fmap_145[15:0]) +
	( 3'sd 3) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 7) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 6) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 3'sd 3) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 3'sd 3) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 3'sd 2) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 3'sd 2) * $signed(input_fmap_203[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 5) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 6) * $signed(input_fmap_232[15:0]) +
	( 3'sd 3) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 2'sd 1) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_241;
assign conv_mac_241 = 
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 5'sd 8) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 7) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 5) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 4'sd 7) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 6) * $signed(input_fmap_55[15:0]) +
	( 3'sd 2) * $signed(input_fmap_56[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 6) * $signed(input_fmap_58[15:0]) +
	( 4'sd 4) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 2'sd 1) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 3) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 3'sd 3) * $signed(input_fmap_90[15:0]) +
	( 2'sd 1) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 7) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 2) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 4'sd 5) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 5'sd 8) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 3'sd 3) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 7) * $signed(input_fmap_136[15:0]) +
	( 4'sd 4) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 5) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 2'sd 1) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 5) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 3'sd 2) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 5) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 7) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 3) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 3'sd 2) * $signed(input_fmap_197[15:0]) +
	( 4'sd 4) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 5'sd 8) * $signed(input_fmap_200[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 6) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 4) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_240[15:0]) +
	( 4'sd 7) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 7) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_242;
assign conv_mac_242 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 4) * $signed(input_fmap_1[15:0]) +
	( 3'sd 2) * $signed(input_fmap_2[15:0]) +
	( 3'sd 3) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 7) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 7) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 7) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 4'sd 5) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 4'sd 7) * $signed(input_fmap_51[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 3'sd 2) * $signed(input_fmap_55[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 5'sd 8) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 5'sd 8) * $signed(input_fmap_83[15:0]) +
	( 4'sd 7) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 4'sd 6) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 5'sd 8) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 5'sd 8) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 3'sd 3) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 5'sd 8) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 4'sd 5) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 7) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 3'sd 3) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 6) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 4'sd 6) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 5'sd 8) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 3'sd 2) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 2'sd 1) * $signed(input_fmap_195[15:0]) +
	( 2'sd 1) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 3) * $signed(input_fmap_203[15:0]) +
	( 3'sd 3) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 5'sd 8) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 6) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 3'sd 3) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_228[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 3'sd 2) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 5) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_238[15:0]) +
	( 4'sd 7) * $signed(input_fmap_239[15:0]) +
	( 3'sd 3) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_243;
assign conv_mac_243 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 5'sd 8) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 4'sd 7) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 2'sd 1) * $signed(input_fmap_20[15:0]) +
	( 5'sd 8) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 4'sd 5) * $signed(input_fmap_32[15:0]) +
	( 4'sd 5) * $signed(input_fmap_33[15:0]) +
	( 4'sd 7) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 4'sd 5) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 4'sd 7) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 5'sd 8) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 4) * $signed(input_fmap_60[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 3'sd 2) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 5'sd 8) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 4) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 6) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 5) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 6) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 4) * $signed(input_fmap_96[15:0]) +
	( 4'sd 6) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 7) * $signed(input_fmap_103[15:0]) +
	( 2'sd 1) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 3'sd 2) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 4'sd 6) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 5'sd 8) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 2'sd 1) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 4'sd 7) * $signed(input_fmap_132[15:0]) +
	( 2'sd 1) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 3'sd 2) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 4'sd 6) * $signed(input_fmap_138[15:0]) +
	( 4'sd 7) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 5) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 5'sd 8) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 3) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 3'sd 2) * $signed(input_fmap_169[15:0]) +
	( 4'sd 5) * $signed(input_fmap_170[15:0]) +
	( 4'sd 7) * $signed(input_fmap_171[15:0]) +
	( 5'sd 8) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 7) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 3'sd 2) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 3'sd 3) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 7) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 5'sd 8) * $signed(input_fmap_206[15:0]) +
	( 4'sd 6) * $signed(input_fmap_207[15:0]) +
	( 2'sd 1) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 5) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 4) * $signed(input_fmap_216[15:0]) +
	( 4'sd 7) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 3) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 3'sd 2) * $signed(input_fmap_227[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 3'sd 2) * $signed(input_fmap_229[15:0]) +
	( 2'sd 1) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 5'sd 8) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_235[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 5'sd 8) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 6) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 7) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_244;
assign conv_mac_244 = 
	( 2'sd 1) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 4'sd 7) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 7) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 3'sd 2) * $signed(input_fmap_20[15:0]) +
	( 4'sd 6) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 3'sd 3) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 4'sd 7) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 5'sd 8) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 3'sd 3) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 6) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 2'sd 1) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 5'sd 8) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 4'sd 5) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 4'sd 5) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 2'sd 1) * $signed(input_fmap_98[15:0]) +
	( 3'sd 3) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_100[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 3'sd 2) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 4) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 2'sd 1) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 2'sd 1) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 4) * $signed(input_fmap_142[15:0]) +
	( 2'sd 1) * $signed(input_fmap_143[15:0]) +
	( 4'sd 6) * $signed(input_fmap_144[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 2'sd 1) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 3'sd 2) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 6) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 4'sd 4) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 4'sd 4) * $signed(input_fmap_184[15:0]) +
	( 4'sd 6) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 3'sd 2) * $signed(input_fmap_187[15:0]) +
	( 2'sd 1) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 4'sd 4) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 4'sd 7) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 3'sd 3) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 5'sd 8) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 4'sd 7) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 4'sd 6) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 2'sd 1) * $signed(input_fmap_232[15:0]) +
	( 4'sd 4) * $signed(input_fmap_233[15:0]) +
	( 4'sd 7) * $signed(input_fmap_234[15:0]) +
	( 4'sd 4) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 6) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 4) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_244[15:0]) +
	( 3'sd 3) * $signed(input_fmap_245[15:0]) +
	( 4'sd 5) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 4) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_245;
assign conv_mac_245 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 3'sd 2) * $signed(input_fmap_1[15:0]) +
	( 4'sd 7) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 5'sd 8) * $signed(input_fmap_9[15:0]) +
	( 4'sd 5) * $signed(input_fmap_10[15:0]) +
	( 2'sd 1) * $signed(input_fmap_11[15:0]) +
	( 3'sd 2) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 5) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 4'sd 7) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 3) * $signed(input_fmap_23[15:0]) +
	( 3'sd 3) * $signed(input_fmap_24[15:0]) +
	( 3'sd 2) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 2'sd 1) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 4'sd 7) * $signed(input_fmap_38[15:0]) +
	( 4'sd 4) * $signed(input_fmap_39[15:0]) +
	( 4'sd 4) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 5) * $signed(input_fmap_42[15:0]) +
	( 5'sd 8) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 2'sd 1) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 6) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_49[15:0]) +
	( 5'sd 8) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 5'sd 8) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 4'sd 7) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 4'sd 7) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_82[15:0]) +
	( 2'sd 1) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 3'sd 2) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 3) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 3'sd 3) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 3'sd 2) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 2'sd 1) * $signed(input_fmap_103[15:0]) +
	( 3'sd 3) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 4'sd 5) * $signed(input_fmap_113[15:0]) +
	( 5'sd 8) * $signed(input_fmap_114[15:0]) +
	( 4'sd 5) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 4'sd 7) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 7) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 2'sd 1) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 5'sd 8) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 4) * $signed(input_fmap_143[15:0]) +
	( 5'sd 8) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 3'sd 3) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 4'sd 5) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 4) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 4) * $signed(input_fmap_156[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 4'sd 7) * $signed(input_fmap_159[15:0]) +
	( 3'sd 2) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 3'sd 3) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 4'sd 6) * $signed(input_fmap_167[15:0]) +
	( 2'sd 1) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 2'sd 1) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 3'sd 3) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 6) * $signed(input_fmap_182[15:0]) +
	( 4'sd 5) * $signed(input_fmap_184[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 6) * $signed(input_fmap_189[15:0]) +
	( 4'sd 7) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 2'sd 1) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 4) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_205[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 5'sd 8) * $signed(input_fmap_210[15:0]) +
	( 3'sd 2) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 4'sd 5) * $signed(input_fmap_216[15:0]) +
	( 5'sd 8) * $signed(input_fmap_217[15:0]) +
	( 4'sd 6) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 4'sd 7) * $signed(input_fmap_222[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 3'sd 2) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 5'sd 8) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 5) * $signed(input_fmap_235[15:0]) +
	( 5'sd 8) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 4'sd 6) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 4'sd 7) * $signed(input_fmap_251[15:0]) +
	( 4'sd 4) * $signed(input_fmap_252[15:0]) +
	( 2'sd 1) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]);

logic signed [31:0] conv_mac_246;
assign conv_mac_246 = 
	( 4'sd 6) * $signed(input_fmap_0[15:0]) +
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 4'sd 6) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 7) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 2) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 4'sd 5) * $signed(input_fmap_14[15:0]) +
	( 3'sd 2) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 4'sd 5) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 5'sd 8) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 2'sd 1) * $signed(input_fmap_43[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 5'sd 8) * $signed(input_fmap_47[15:0]) +
	( 2'sd 1) * $signed(input_fmap_48[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 4'sd 4) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 2) * $signed(input_fmap_52[15:0]) +
	( 4'sd 7) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 2'sd 1) * $signed(input_fmap_56[15:0]) +
	( 4'sd 5) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 4'sd 6) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 3'sd 3) * $signed(input_fmap_70[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 2'sd 1) * $signed(input_fmap_73[15:0]) +
	( 5'sd 8) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_77[15:0]) +
	( 4'sd 6) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 5) * $signed(input_fmap_87[15:0]) +
	( 4'sd 4) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 6) * $signed(input_fmap_90[15:0]) +
	( 3'sd 3) * $signed(input_fmap_91[15:0]) +
	( 3'sd 2) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 5'sd 8) * $signed(input_fmap_94[15:0]) +
	( 4'sd 4) * $signed(input_fmap_95[15:0]) +
	( 2'sd 1) * $signed(input_fmap_96[15:0]) +
	( 4'sd 4) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 3'sd 2) * $signed(input_fmap_104[15:0]) +
	( 5'sd 8) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 5'sd 8) * $signed(input_fmap_113[15:0]) +
	( 4'sd 7) * $signed(input_fmap_114[15:0]) +
	( 3'sd 3) * $signed(input_fmap_115[15:0]) +
	( 4'sd 6) * $signed(input_fmap_116[15:0]) +
	( 3'sd 3) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 2) * $signed(input_fmap_119[15:0]) +
	( 4'sd 7) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 3'sd 3) * $signed(input_fmap_125[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 2'sd 1) * $signed(input_fmap_131[15:0]) +
	( 5'sd 8) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 4'sd 6) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 4'sd 5) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_145[15:0]) +
	( 4'sd 4) * $signed(input_fmap_146[15:0]) +
	( 3'sd 2) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 2'sd 1) * $signed(input_fmap_151[15:0]) +
	( 4'sd 4) * $signed(input_fmap_152[15:0]) +
	( 4'sd 5) * $signed(input_fmap_153[15:0]) +
	( 4'sd 5) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 3'sd 3) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 4'sd 6) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 4) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 2'sd 1) * $signed(input_fmap_171[15:0]) +
	( 3'sd 3) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 6) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 6) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 3'sd 2) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 4'sd 6) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 4'sd 5) * $signed(input_fmap_198[15:0]) +
	( 4'sd 7) * $signed(input_fmap_199[15:0]) +
	( 3'sd 2) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 5'sd 8) * $signed(input_fmap_204[15:0]) +
	( 3'sd 3) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 7) * $signed(input_fmap_209[15:0]) +
	( 3'sd 3) * $signed(input_fmap_210[15:0]) +
	( 3'sd 3) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 5'sd 8) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 4'sd 4) * $signed(input_fmap_223[15:0]) +
	( 4'sd 6) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 6) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 5) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 2'sd 1) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 4'sd 7) * $signed(input_fmap_247[15:0]) +
	( 4'sd 5) * $signed(input_fmap_248[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_254[15:0]) +
	( 4'sd 6) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_247;
assign conv_mac_247 = 
	( 3'sd 3) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 4) * $signed(input_fmap_3[15:0]) +
	( 4'sd 5) * $signed(input_fmap_4[15:0]) +
	( 3'sd 2) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 5) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_13[15:0]) +
	( 3'sd 3) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 4'sd 6) * $signed(input_fmap_19[15:0]) +
	( 4'sd 7) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 3'sd 2) * $signed(input_fmap_23[15:0]) +
	( 4'sd 6) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 7) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_35[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 5) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_41[15:0]) +
	( 4'sd 7) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 7) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 2'sd 1) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_52[15:0]) +
	( 3'sd 2) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 5'sd 8) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 2) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 3'sd 2) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 3'sd 2) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 5'sd 8) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 4'sd 4) * $signed(input_fmap_78[15:0]) +
	( 4'sd 6) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 6) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 4'sd 5) * $signed(input_fmap_90[15:0]) +
	( 3'sd 2) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_98[15:0]) +
	( 4'sd 6) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 7) * $signed(input_fmap_106[15:0]) +
	( 4'sd 7) * $signed(input_fmap_107[15:0]) +
	( 4'sd 6) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 7) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 3'sd 3) * $signed(input_fmap_119[15:0]) +
	( 4'sd 6) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 3) * $signed(input_fmap_123[15:0]) +
	( 5'sd 8) * $signed(input_fmap_124[15:0]) +
	( 3'sd 2) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 6) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 7) * $signed(input_fmap_138[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 4'sd 7) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 4'sd 6) * $signed(input_fmap_148[15:0]) +
	( 2'sd 1) * $signed(input_fmap_149[15:0]) +
	( 4'sd 7) * $signed(input_fmap_150[15:0]) +
	( 3'sd 3) * $signed(input_fmap_151[15:0]) +
	( 3'sd 3) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 2'sd 1) * $signed(input_fmap_155[15:0]) +
	( 3'sd 3) * $signed(input_fmap_156[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 5) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 2'sd 1) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 3'sd 3) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 3'sd 2) * $signed(input_fmap_182[15:0]) +
	( 5'sd 8) * $signed(input_fmap_183[15:0]) +
	( 3'sd 2) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 5'sd 8) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 2'sd 1) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_204[15:0]) +
	( 4'sd 4) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 4'sd 7) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 6) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 5'sd 8) * $signed(input_fmap_230[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 2'sd 1) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 2'sd 1) * $signed(input_fmap_238[15:0]) +
	( 4'sd 4) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 7) * $signed(input_fmap_246[15:0]) +
	( 4'sd 5) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 3'sd 3) * $signed(input_fmap_250[15:0]) +
	( 4'sd 6) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_248;
assign conv_mac_248 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 3'sd 2) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 3'sd 3) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 4'sd 6) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 5) * $signed(input_fmap_12[15:0]) +
	( 4'sd 6) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 3'sd 2) * $signed(input_fmap_16[15:0]) +
	( 3'sd 2) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 4'sd 5) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 5'sd 8) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 4) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 3'sd 3) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 2) * $signed(input_fmap_32[15:0]) +
	( 4'sd 7) * $signed(input_fmap_33[15:0]) +
	( 3'sd 2) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 5) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 2'sd 1) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 4'sd 5) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 2'sd 1) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 7) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 3'sd 3) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 4'sd 5) * $signed(input_fmap_65[15:0]) +
	( 3'sd 2) * $signed(input_fmap_66[15:0]) +
	( 4'sd 6) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 7) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_71[15:0]) +
	( 4'sd 7) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 4'sd 4) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 4'sd 4) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 2'sd 1) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 7) * $signed(input_fmap_80[15:0]) +
	( 3'sd 2) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_85[15:0]) +
	( 4'sd 6) * $signed(input_fmap_86[15:0]) +
	( 4'sd 7) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 4) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 4) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 4'sd 7) * $signed(input_fmap_101[15:0]) +
	( 5'sd 8) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 5) * $signed(input_fmap_105[15:0]) +
	( 3'sd 2) * $signed(input_fmap_106[15:0]) +
	( 3'sd 3) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 4'sd 7) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 3'sd 3) * $signed(input_fmap_112[15:0]) +
	( 3'sd 3) * $signed(input_fmap_113[15:0]) +
	( 3'sd 3) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 2'sd 1) * $signed(input_fmap_122[15:0]) +
	( 3'sd 2) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 3'sd 2) * $signed(input_fmap_132[15:0]) +
	( 4'sd 5) * $signed(input_fmap_133[15:0]) +
	( 3'sd 2) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 3'sd 3) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 5'sd 8) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 4'sd 6) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 3'sd 2) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 5'sd 8) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 7) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 5'sd 8) * $signed(input_fmap_165[15:0]) +
	( 2'sd 1) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 4'sd 5) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_175[15:0]) +
	( 3'sd 3) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 4'sd 7) * $signed(input_fmap_180[15:0]) +
	( 5'sd 8) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 4'sd 5) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 4'sd 5) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 3'sd 3) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 4'sd 4) * $signed(input_fmap_196[15:0]) +
	( 3'sd 3) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_199[15:0]) +
	( 2'sd 1) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 4) * $signed(input_fmap_202[15:0]) +
	( 4'sd 7) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 3'sd 2) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 2'sd 1) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 2'sd 1) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 4'sd 6) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 5) * $signed(input_fmap_224[15:0]) +
	( 2'sd 1) * $signed(input_fmap_225[15:0]) +
	( 5'sd 8) * $signed(input_fmap_227[15:0]) +
	( 4'sd 4) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 2) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 3'sd 2) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 4'sd 5) * $signed(input_fmap_237[15:0]) +
	( 4'sd 4) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 7) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 4'sd 7) * $signed(input_fmap_244[15:0]) +
	( 4'sd 5) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 5) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 4'sd 5) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 5'sd 8) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_249;
assign conv_mac_249 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 4'sd 5) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_3[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 4'sd 4) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_13[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 4) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 4'sd 4) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 4'sd 4) * $signed(input_fmap_21[15:0]) +
	( 4'sd 5) * $signed(input_fmap_22[15:0]) +
	( 4'sd 7) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 3) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 3'sd 2) * $signed(input_fmap_33[15:0]) +
	( 4'sd 6) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 3'sd 3) * $signed(input_fmap_37[15:0]) +
	( 2'sd 1) * $signed(input_fmap_38[15:0]) +
	( 4'sd 5) * $signed(input_fmap_39[15:0]) +
	( 4'sd 5) * $signed(input_fmap_40[15:0]) +
	( 4'sd 4) * $signed(input_fmap_41[15:0]) +
	( 3'sd 2) * $signed(input_fmap_42[15:0]) +
	( 4'sd 5) * $signed(input_fmap_43[15:0]) +
	( 4'sd 6) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 4'sd 4) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 3'sd 2) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 5) * $signed(input_fmap_58[15:0]) +
	( 5'sd 8) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_60[15:0]) +
	( 4'sd 7) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 3'sd 3) * $signed(input_fmap_63[15:0]) +
	( 4'sd 6) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 6) * $signed(input_fmap_66[15:0]) +
	( 5'sd 8) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 6) * $signed(input_fmap_69[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 3'sd 3) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 4'sd 7) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 2'sd 1) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 5'sd 8) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 3'sd 2) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 4) * $signed(input_fmap_86[15:0]) +
	( 4'sd 6) * $signed(input_fmap_87[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 4'sd 6) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 2'sd 1) * $signed(input_fmap_94[15:0]) +
	( 3'sd 2) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 2) * $signed(input_fmap_97[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 5) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 3'sd 3) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 3'sd 3) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 3'sd 2) * $signed(input_fmap_113[15:0]) +
	( 2'sd 1) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 3'sd 2) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 4'sd 5) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_122[15:0]) +
	( 4'sd 4) * $signed(input_fmap_123[15:0]) +
	( 4'sd 4) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 2) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 2'sd 1) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 5'sd 8) * $signed(input_fmap_140[15:0]) +
	( 4'sd 7) * $signed(input_fmap_141[15:0]) +
	( 3'sd 3) * $signed(input_fmap_142[15:0]) +
	( 4'sd 6) * $signed(input_fmap_143[15:0]) +
	( 4'sd 7) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_146[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 4'sd 7) * $signed(input_fmap_148[15:0]) +
	( 3'sd 3) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 4'sd 5) * $signed(input_fmap_152[15:0]) +
	( 2'sd 1) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 7) * $signed(input_fmap_155[15:0]) +
	( 4'sd 6) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 4'sd 5) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 5) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 4'sd 4) * $signed(input_fmap_164[15:0]) +
	( 4'sd 6) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 7) * $signed(input_fmap_172[15:0]) +
	( 5'sd 8) * $signed(input_fmap_173[15:0]) +
	( 5'sd 8) * $signed(input_fmap_174[15:0]) +
	( 4'sd 6) * $signed(input_fmap_175[15:0]) +
	( 3'sd 2) * $signed(input_fmap_176[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 5'sd 8) * $signed(input_fmap_178[15:0]) +
	( 4'sd 7) * $signed(input_fmap_179[15:0]) +
	( 3'sd 3) * $signed(input_fmap_180[15:0]) +
	( 4'sd 7) * $signed(input_fmap_181[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 4'sd 6) * $signed(input_fmap_187[15:0]) +
	( 5'sd 8) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 4'sd 7) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 2'sd 1) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 6) * $signed(input_fmap_195[15:0]) +
	( 5'sd 8) * $signed(input_fmap_196[15:0]) +
	( 2'sd 1) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 4'sd 7) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_205[15:0]) +
	( 3'sd 3) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 5) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 4) * $signed(input_fmap_215[15:0]) +
	( 4'sd 6) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 5) * $signed(input_fmap_220[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 2'sd 1) * $signed(input_fmap_223[15:0]) +
	( 5'sd 8) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 4'sd 7) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_228[15:0]) +
	( 4'sd 4) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 3'sd 3) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 2) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_237[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 3'sd 3) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 4) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 5'sd 8) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 3'sd 3) * $signed(input_fmap_252[15:0]) +
	( 4'sd 7) * $signed(input_fmap_253[15:0]) +
	( 4'sd 4) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_250;
assign conv_mac_250 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 7) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 3) * $signed(input_fmap_7[15:0]) +
	( 4'sd 4) * $signed(input_fmap_9[15:0]) +
	( 5'sd 8) * $signed(input_fmap_10[15:0]) +
	( 4'sd 4) * $signed(input_fmap_11[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 5'sd 8) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 5) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 4) * $signed(input_fmap_23[15:0]) +
	( 3'sd 2) * $signed(input_fmap_24[15:0]) +
	( 4'sd 6) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 7) * $signed(input_fmap_27[15:0]) +
	( 3'sd 3) * $signed(input_fmap_28[15:0]) +
	( 2'sd 1) * $signed(input_fmap_29[15:0]) +
	( 5'sd 8) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 4'sd 4) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 4'sd 4) * $signed(input_fmap_35[15:0]) +
	( 4'sd 7) * $signed(input_fmap_36[15:0]) +
	( 2'sd 1) * $signed(input_fmap_37[15:0]) +
	( 4'sd 4) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_42[15:0]) +
	( 4'sd 4) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 4'sd 7) * $signed(input_fmap_47[15:0]) +
	( 4'sd 7) * $signed(input_fmap_48[15:0]) +
	( 4'sd 4) * $signed(input_fmap_49[15:0]) +
	( 3'sd 3) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 3'sd 3) * $signed(input_fmap_52[15:0]) +
	( 3'sd 3) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 5'sd 8) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 3'sd 3) * $signed(input_fmap_60[15:0]) +
	( 4'sd 4) * $signed(input_fmap_61[15:0]) +
	( 2'sd 1) * $signed(input_fmap_63[15:0]) +
	( 2'sd 1) * $signed(input_fmap_64[15:0]) +
	( 5'sd 8) * $signed(input_fmap_65[15:0]) +
	( 3'sd 3) * $signed(input_fmap_66[15:0]) +
	( 4'sd 4) * $signed(input_fmap_67[15:0]) +
	( 4'sd 7) * $signed(input_fmap_68[15:0]) +
	( 2'sd 1) * $signed(input_fmap_69[15:0]) +
	( 2'sd 1) * $signed(input_fmap_70[15:0]) +
	( 4'sd 7) * $signed(input_fmap_71[15:0]) +
	( 4'sd 4) * $signed(input_fmap_72[15:0]) +
	( 4'sd 6) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 3'sd 3) * $signed(input_fmap_76[15:0]) +
	( 4'sd 6) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 2'sd 1) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 3'sd 3) * $signed(input_fmap_84[15:0]) +
	( 2'sd 1) * $signed(input_fmap_85[15:0]) +
	( 4'sd 7) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 5'sd 8) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_98[15:0]) +
	( 2'sd 1) * $signed(input_fmap_100[15:0]) +
	( 3'sd 3) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_106[15:0]) +
	( 2'sd 1) * $signed(input_fmap_107[15:0]) +
	( 3'sd 3) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 2'sd 1) * $signed(input_fmap_110[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 5'sd 8) * $signed(input_fmap_115[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_117[15:0]) +
	( 2'sd 1) * $signed(input_fmap_118[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 4'sd 7) * $signed(input_fmap_129[15:0]) +
	( 4'sd 5) * $signed(input_fmap_130[15:0]) +
	( 4'sd 6) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 6) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 4) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 4) * $signed(input_fmap_140[15:0]) +
	( 4'sd 6) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 3) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 3'sd 2) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 6) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 5) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 4) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 4'sd 6) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 3'sd 3) * $signed(input_fmap_160[15:0]) +
	( 2'sd 1) * $signed(input_fmap_161[15:0]) +
	( 4'sd 4) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 5) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 3'sd 2) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_168[15:0]) +
	( 4'sd 4) * $signed(input_fmap_169[15:0]) +
	( 5'sd 8) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 4'sd 6) * $signed(input_fmap_172[15:0]) +
	( 4'sd 5) * $signed(input_fmap_173[15:0]) +
	( 3'sd 2) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 5) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_177[15:0]) +
	( 3'sd 2) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 5) * $signed(input_fmap_180[15:0]) +
	( 4'sd 6) * $signed(input_fmap_181[15:0]) +
	( 5'sd 8) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 5'sd 8) * $signed(input_fmap_185[15:0]) +
	( 5'sd 8) * $signed(input_fmap_186[15:0]) +
	( 4'sd 7) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 3'sd 3) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 5'sd 8) * $signed(input_fmap_194[15:0]) +
	( 3'sd 2) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 5'sd 8) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 5'sd 8) * $signed(input_fmap_201[15:0]) +
	( 4'sd 5) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 6) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 7) * $signed(input_fmap_207[15:0]) +
	( 4'sd 6) * $signed(input_fmap_208[15:0]) +
	( 4'sd 5) * $signed(input_fmap_209[15:0]) +
	( 2'sd 1) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 4'sd 6) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 4'sd 5) * $signed(input_fmap_218[15:0]) +
	( 4'sd 7) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 4'sd 7) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 4'sd 5) * $signed(input_fmap_227[15:0]) +
	( 4'sd 6) * $signed(input_fmap_229[15:0]) +
	( 4'sd 6) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 6) * $signed(input_fmap_236[15:0]) +
	( 2'sd 1) * $signed(input_fmap_237[15:0]) +
	( 5'sd 8) * $signed(input_fmap_238[15:0]) +
	( 3'sd 3) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 2'sd 1) * $signed(input_fmap_242[15:0]) +
	( 3'sd 2) * $signed(input_fmap_243[15:0]) +
	( 2'sd 1) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 3'sd 2) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_248[15:0]) +
	( 3'sd 2) * $signed(input_fmap_249[15:0]) +
	( 4'sd 7) * $signed(input_fmap_250[15:0]) +
	( 4'sd 4) * $signed(input_fmap_251[15:0]) +
	( 4'sd 7) * $signed(input_fmap_252[15:0]) +
	( 4'sd 5) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_251;
assign conv_mac_251 = 
	( 4'sd 7) * $signed(input_fmap_0[15:0]) +
	( 2'sd 1) * $signed(input_fmap_1[15:0]) +
	( 5'sd 8) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 4'sd 5) * $signed(input_fmap_7[15:0]) +
	( 4'sd 5) * $signed(input_fmap_8[15:0]) +
	( 4'sd 7) * $signed(input_fmap_9[15:0]) +
	( 4'sd 4) * $signed(input_fmap_10[15:0]) +
	( 4'sd 5) * $signed(input_fmap_11[15:0]) +
	( 4'sd 6) * $signed(input_fmap_12[15:0]) +
	( 4'sd 7) * $signed(input_fmap_13[15:0]) +
	( 2'sd 1) * $signed(input_fmap_14[15:0]) +
	( 4'sd 7) * $signed(input_fmap_15[15:0]) +
	( 2'sd 1) * $signed(input_fmap_16[15:0]) +
	( 3'sd 3) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 5) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 4'sd 5) * $signed(input_fmap_24[15:0]) +
	( 5'sd 8) * $signed(input_fmap_25[15:0]) +
	( 4'sd 7) * $signed(input_fmap_26[15:0]) +
	( 4'sd 5) * $signed(input_fmap_27[15:0]) +
	( 4'sd 7) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 5) * $signed(input_fmap_30[15:0]) +
	( 3'sd 3) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 5'sd 8) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 3'sd 2) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 3'sd 2) * $signed(input_fmap_38[15:0]) +
	( 4'sd 6) * $signed(input_fmap_39[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 2'sd 1) * $signed(input_fmap_44[15:0]) +
	( 4'sd 5) * $signed(input_fmap_45[15:0]) +
	( 4'sd 4) * $signed(input_fmap_46[15:0]) +
	( 2'sd 1) * $signed(input_fmap_47[15:0]) +
	( 4'sd 5) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 3'sd 3) * $signed(input_fmap_51[15:0]) +
	( 5'sd 8) * $signed(input_fmap_52[15:0]) +
	( 4'sd 6) * $signed(input_fmap_53[15:0]) +
	( 3'sd 3) * $signed(input_fmap_54[15:0]) +
	( 4'sd 4) * $signed(input_fmap_56[15:0]) +
	( 3'sd 2) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 3'sd 2) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 2) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 3'sd 3) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 4'sd 5) * $signed(input_fmap_67[15:0]) +
	( 4'sd 6) * $signed(input_fmap_68[15:0]) +
	( 5'sd 8) * $signed(input_fmap_69[15:0]) +
	( 3'sd 2) * $signed(input_fmap_70[15:0]) +
	( 4'sd 4) * $signed(input_fmap_71[15:0]) +
	( 3'sd 3) * $signed(input_fmap_72[15:0]) +
	( 4'sd 5) * $signed(input_fmap_73[15:0]) +
	( 4'sd 5) * $signed(input_fmap_74[15:0]) +
	( 4'sd 6) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 5) * $signed(input_fmap_77[15:0]) +
	( 4'sd 5) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 4'sd 7) * $signed(input_fmap_83[15:0]) +
	( 3'sd 2) * $signed(input_fmap_84[15:0]) +
	( 3'sd 3) * $signed(input_fmap_85[15:0]) +
	( 5'sd 8) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 3'sd 3) * $signed(input_fmap_88[15:0]) +
	( 4'sd 5) * $signed(input_fmap_89[15:0]) +
	( 4'sd 7) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 5'sd 8) * $signed(input_fmap_92[15:0]) +
	( 4'sd 5) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 4'sd 5) * $signed(input_fmap_95[15:0]) +
	( 3'sd 2) * $signed(input_fmap_96[15:0]) +
	( 4'sd 5) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 4'sd 5) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 5'sd 8) * $signed(input_fmap_101[15:0]) +
	( 4'sd 7) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 7) * $signed(input_fmap_110[15:0]) +
	( 4'sd 5) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 6) * $signed(input_fmap_115[15:0]) +
	( 4'sd 5) * $signed(input_fmap_116[15:0]) +
	( 5'sd 8) * $signed(input_fmap_118[15:0]) +
	( 2'sd 1) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 6) * $signed(input_fmap_124[15:0]) +
	( 4'sd 5) * $signed(input_fmap_125[15:0]) +
	( 2'sd 1) * $signed(input_fmap_126[15:0]) +
	( 4'sd 5) * $signed(input_fmap_127[15:0]) +
	( 2'sd 1) * $signed(input_fmap_128[15:0]) +
	( 3'sd 2) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 5) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 7) * $signed(input_fmap_133[15:0]) +
	( 4'sd 7) * $signed(input_fmap_134[15:0]) +
	( 4'sd 6) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 6) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 3'sd 2) * $signed(input_fmap_141[15:0]) +
	( 3'sd 2) * $signed(input_fmap_142[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 5) * $signed(input_fmap_145[15:0]) +
	( 4'sd 5) * $signed(input_fmap_147[15:0]) +
	( 2'sd 1) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 6) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 3'sd 3) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 7) * $signed(input_fmap_156[15:0]) +
	( 3'sd 2) * $signed(input_fmap_157[15:0]) +
	( 3'sd 2) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 3'sd 2) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 3'sd 2) * $signed(input_fmap_165[15:0]) +
	( 4'sd 7) * $signed(input_fmap_166[15:0]) +
	( 4'sd 7) * $signed(input_fmap_167[15:0]) +
	( 4'sd 6) * $signed(input_fmap_168[15:0]) +
	( 4'sd 5) * $signed(input_fmap_169[15:0]) +
	( 3'sd 2) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 3'sd 3) * $signed(input_fmap_174[15:0]) +
	( 2'sd 1) * $signed(input_fmap_175[15:0]) +
	( 4'sd 4) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 5) * $signed(input_fmap_179[15:0]) +
	( 4'sd 4) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 4) * $signed(input_fmap_185[15:0]) +
	( 3'sd 2) * $signed(input_fmap_186[15:0]) +
	( 4'sd 5) * $signed(input_fmap_187[15:0]) +
	( 3'sd 3) * $signed(input_fmap_188[15:0]) +
	( 4'sd 5) * $signed(input_fmap_189[15:0]) +
	( 3'sd 2) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 4'sd 7) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 4'sd 7) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 6) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 2'sd 1) * $signed(input_fmap_204[15:0]) +
	( 5'sd 8) * $signed(input_fmap_205[15:0]) +
	( 4'sd 6) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 3'sd 2) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_209[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 2'sd 1) * $signed(input_fmap_213[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_217[15:0]) +
	( 5'sd 8) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 4'sd 7) * $signed(input_fmap_220[15:0]) +
	( 3'sd 3) * $signed(input_fmap_221[15:0]) +
	( 2'sd 1) * $signed(input_fmap_222[15:0]) +
	( 4'sd 5) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 5) * $signed(input_fmap_225[15:0]) +
	( 3'sd 3) * $signed(input_fmap_226[15:0]) +
	( 4'sd 7) * $signed(input_fmap_227[15:0]) +
	( 4'sd 7) * $signed(input_fmap_228[15:0]) +
	( 4'sd 7) * $signed(input_fmap_229[15:0]) +
	( 4'sd 7) * $signed(input_fmap_230[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 5'sd 8) * $signed(input_fmap_233[15:0]) +
	( 2'sd 1) * $signed(input_fmap_234[15:0]) +
	( 2'sd 1) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 5) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 3'sd 3) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 4) * $signed(input_fmap_245[15:0]) +
	( 3'sd 3) * $signed(input_fmap_246[15:0]) +
	( 2'sd 1) * $signed(input_fmap_247[15:0]) +
	( 4'sd 7) * $signed(input_fmap_248[15:0]) +
	( 2'sd 1) * $signed(input_fmap_249[15:0]) +
	( 4'sd 6) * $signed(input_fmap_250[15:0]) +
	( 3'sd 3) * $signed(input_fmap_251[15:0]) +
	( 3'sd 2) * $signed(input_fmap_252[15:0]) +
	( 3'sd 2) * $signed(input_fmap_253[15:0]) +
	( 3'sd 3) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_252;
assign conv_mac_252 = 
	( 4'sd 5) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 2'sd 1) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 4) * $signed(input_fmap_5[15:0]) +
	( 2'sd 1) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 2'sd 1) * $signed(input_fmap_9[15:0]) +
	( 3'sd 2) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 2'sd 1) * $signed(input_fmap_12[15:0]) +
	( 4'sd 4) * $signed(input_fmap_13[15:0]) +
	( 4'sd 4) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_15[15:0]) +
	( 3'sd 3) * $signed(input_fmap_16[15:0]) +
	( 2'sd 1) * $signed(input_fmap_17[15:0]) +
	( 3'sd 2) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 3'sd 3) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 4) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 5) * $signed(input_fmap_28[15:0]) +
	( 4'sd 4) * $signed(input_fmap_29[15:0]) +
	( 4'sd 7) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 4'sd 6) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 4'sd 5) * $signed(input_fmap_36[15:0]) +
	( 4'sd 7) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_39[15:0]) +
	( 2'sd 1) * $signed(input_fmap_40[15:0]) +
	( 3'sd 3) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 6) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 6) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 3'sd 3) * $signed(input_fmap_47[15:0]) +
	( 3'sd 3) * $signed(input_fmap_48[15:0]) +
	( 4'sd 6) * $signed(input_fmap_49[15:0]) +
	( 4'sd 6) * $signed(input_fmap_50[15:0]) +
	( 3'sd 2) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 7) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 4'sd 4) * $signed(input_fmap_57[15:0]) +
	( 4'sd 7) * $signed(input_fmap_58[15:0]) +
	( 4'sd 6) * $signed(input_fmap_59[15:0]) +
	( 4'sd 7) * $signed(input_fmap_60[15:0]) +
	( 3'sd 3) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 3'sd 2) * $signed(input_fmap_63[15:0]) +
	( 4'sd 7) * $signed(input_fmap_64[15:0]) +
	( 3'sd 3) * $signed(input_fmap_65[15:0]) +
	( 5'sd 8) * $signed(input_fmap_66[15:0]) +
	( 3'sd 2) * $signed(input_fmap_67[15:0]) +
	( 4'sd 4) * $signed(input_fmap_68[15:0]) +
	( 4'sd 5) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_71[15:0]) +
	( 4'sd 6) * $signed(input_fmap_72[15:0]) +
	( 3'sd 2) * $signed(input_fmap_73[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 5'sd 8) * $signed(input_fmap_76[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 4) * $signed(input_fmap_79[15:0]) +
	( 2'sd 1) * $signed(input_fmap_80[15:0]) +
	( 4'sd 7) * $signed(input_fmap_81[15:0]) +
	( 4'sd 6) * $signed(input_fmap_82[15:0]) +
	( 4'sd 4) * $signed(input_fmap_83[15:0]) +
	( 4'sd 6) * $signed(input_fmap_84[15:0]) +
	( 4'sd 6) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 4'sd 5) * $signed(input_fmap_88[15:0]) +
	( 3'sd 2) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 4'sd 7) * $signed(input_fmap_92[15:0]) +
	( 4'sd 6) * $signed(input_fmap_93[15:0]) +
	( 3'sd 3) * $signed(input_fmap_94[15:0]) +
	( 5'sd 8) * $signed(input_fmap_95[15:0]) +
	( 4'sd 5) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 4'sd 7) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 4) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 5) * $signed(input_fmap_104[15:0]) +
	( 4'sd 7) * $signed(input_fmap_105[15:0]) +
	( 4'sd 4) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 5) * $signed(input_fmap_108[15:0]) +
	( 4'sd 5) * $signed(input_fmap_109[15:0]) +
	( 4'sd 5) * $signed(input_fmap_110[15:0]) +
	( 4'sd 7) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 3'sd 2) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 6) * $signed(input_fmap_117[15:0]) +
	( 4'sd 4) * $signed(input_fmap_118[15:0]) +
	( 5'sd 8) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 3'sd 2) * $signed(input_fmap_121[15:0]) +
	( 4'sd 6) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 4'sd 5) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 4'sd 6) * $signed(input_fmap_127[15:0]) +
	( 4'sd 6) * $signed(input_fmap_128[15:0]) +
	( 4'sd 6) * $signed(input_fmap_129[15:0]) +
	( 3'sd 2) * $signed(input_fmap_131[15:0]) +
	( 3'sd 3) * $signed(input_fmap_133[15:0]) +
	( 4'sd 5) * $signed(input_fmap_134[15:0]) +
	( 4'sd 5) * $signed(input_fmap_135[15:0]) +
	( 5'sd 8) * $signed(input_fmap_136[15:0]) +
	( 3'sd 2) * $signed(input_fmap_137[15:0]) +
	( 4'sd 5) * $signed(input_fmap_138[15:0]) +
	( 3'sd 3) * $signed(input_fmap_139[15:0]) +
	( 2'sd 1) * $signed(input_fmap_140[15:0]) +
	( 5'sd 8) * $signed(input_fmap_141[15:0]) +
	( 2'sd 1) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 4'sd 4) * $signed(input_fmap_144[15:0]) +
	( 4'sd 4) * $signed(input_fmap_145[15:0]) +
	( 5'sd 8) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 5) * $signed(input_fmap_151[15:0]) +
	( 4'sd 6) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 3'sd 3) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_155[15:0]) +
	( 2'sd 1) * $signed(input_fmap_156[15:0]) +
	( 2'sd 1) * $signed(input_fmap_157[15:0]) +
	( 4'sd 5) * $signed(input_fmap_158[15:0]) +
	( 2'sd 1) * $signed(input_fmap_159[15:0]) +
	( 2'sd 1) * $signed(input_fmap_160[15:0]) +
	( 4'sd 7) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 2'sd 1) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 4'sd 4) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_167[15:0]) +
	( 3'sd 3) * $signed(input_fmap_168[15:0]) +
	( 3'sd 3) * $signed(input_fmap_169[15:0]) +
	( 2'sd 1) * $signed(input_fmap_170[15:0]) +
	( 3'sd 2) * $signed(input_fmap_171[15:0]) +
	( 3'sd 2) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 3'sd 2) * $signed(input_fmap_177[15:0]) +
	( 4'sd 7) * $signed(input_fmap_178[15:0]) +
	( 4'sd 6) * $signed(input_fmap_180[15:0]) +
	( 3'sd 3) * $signed(input_fmap_181[15:0]) +
	( 2'sd 1) * $signed(input_fmap_182[15:0]) +
	( 4'sd 6) * $signed(input_fmap_183[15:0]) +
	( 3'sd 3) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 4) * $signed(input_fmap_186[15:0]) +
	( 5'sd 8) * $signed(input_fmap_187[15:0]) +
	( 4'sd 7) * $signed(input_fmap_188[15:0]) +
	( 2'sd 1) * $signed(input_fmap_189[15:0]) +
	( 4'sd 6) * $signed(input_fmap_190[15:0]) +
	( 3'sd 2) * $signed(input_fmap_191[15:0]) +
	( 3'sd 3) * $signed(input_fmap_192[15:0]) +
	( 3'sd 3) * $signed(input_fmap_193[15:0]) +
	( 3'sd 2) * $signed(input_fmap_194[15:0]) +
	( 3'sd 3) * $signed(input_fmap_195[15:0]) +
	( 3'sd 2) * $signed(input_fmap_196[15:0]) +
	( 4'sd 6) * $signed(input_fmap_197[15:0]) +
	( 5'sd 8) * $signed(input_fmap_198[15:0]) +
	( 3'sd 2) * $signed(input_fmap_200[15:0]) +
	( 4'sd 5) * $signed(input_fmap_201[15:0]) +
	( 4'sd 7) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 2'sd 1) * $signed(input_fmap_207[15:0]) +
	( 4'sd 4) * $signed(input_fmap_209[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 4'sd 4) * $signed(input_fmap_211[15:0]) +
	( 4'sd 5) * $signed(input_fmap_212[15:0]) +
	( 3'sd 3) * $signed(input_fmap_213[15:0]) +
	( 4'sd 7) * $signed(input_fmap_214[15:0]) +
	( 3'sd 3) * $signed(input_fmap_215[15:0]) +
	( 3'sd 3) * $signed(input_fmap_216[15:0]) +
	( 4'sd 5) * $signed(input_fmap_217[15:0]) +
	( 3'sd 2) * $signed(input_fmap_218[15:0]) +
	( 3'sd 2) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 3'sd 2) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_223[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 5) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 3'sd 3) * $signed(input_fmap_229[15:0]) +
	( 4'sd 4) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 4) * $signed(input_fmap_232[15:0]) +
	( 4'sd 7) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 4'sd 5) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 5) * $signed(input_fmap_240[15:0]) +
	( 3'sd 3) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 6) * $signed(input_fmap_247[15:0]) +
	( 3'sd 3) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 4'sd 5) * $signed(input_fmap_251[15:0]) +
	( 2'sd 1) * $signed(input_fmap_252[15:0]) +
	( 4'sd 6) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 4'sd 5) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_253;
assign conv_mac_253 = 
	( 4'sd 4) * $signed(input_fmap_0[15:0]) +
	( 4'sd 7) * $signed(input_fmap_1[15:0]) +
	( 4'sd 6) * $signed(input_fmap_2[15:0]) +
	( 4'sd 7) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 3'sd 2) * $signed(input_fmap_6[15:0]) +
	( 3'sd 2) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 3) * $signed(input_fmap_9[15:0]) +
	( 4'sd 6) * $signed(input_fmap_10[15:0]) +
	( 5'sd 8) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 4'sd 5) * $signed(input_fmap_15[15:0]) +
	( 4'sd 4) * $signed(input_fmap_16[15:0]) +
	( 4'sd 6) * $signed(input_fmap_17[15:0]) +
	( 4'sd 4) * $signed(input_fmap_18[15:0]) +
	( 3'sd 2) * $signed(input_fmap_19[15:0]) +
	( 4'sd 4) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 6) * $signed(input_fmap_22[15:0]) +
	( 4'sd 6) * $signed(input_fmap_23[15:0]) +
	( 2'sd 1) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 4'sd 4) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 3'sd 2) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 3'sd 3) * $signed(input_fmap_34[15:0]) +
	( 3'sd 3) * $signed(input_fmap_35[15:0]) +
	( 3'sd 3) * $signed(input_fmap_36[15:0]) +
	( 3'sd 2) * $signed(input_fmap_37[15:0]) +
	( 5'sd 8) * $signed(input_fmap_38[15:0]) +
	( 3'sd 3) * $signed(input_fmap_40[15:0]) +
	( 4'sd 7) * $signed(input_fmap_41[15:0]) +
	( 3'sd 3) * $signed(input_fmap_42[15:0]) +
	( 3'sd 3) * $signed(input_fmap_44[15:0]) +
	( 3'sd 3) * $signed(input_fmap_45[15:0]) +
	( 4'sd 6) * $signed(input_fmap_46[15:0]) +
	( 4'sd 4) * $signed(input_fmap_47[15:0]) +
	( 4'sd 4) * $signed(input_fmap_48[15:0]) +
	( 4'sd 7) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 5'sd 8) * $signed(input_fmap_51[15:0]) +
	( 4'sd 6) * $signed(input_fmap_52[15:0]) +
	( 4'sd 5) * $signed(input_fmap_53[15:0]) +
	( 4'sd 6) * $signed(input_fmap_54[15:0]) +
	( 4'sd 5) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 4'sd 6) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 7) * $signed(input_fmap_59[15:0]) +
	( 4'sd 5) * $signed(input_fmap_61[15:0]) +
	( 3'sd 3) * $signed(input_fmap_62[15:0]) +
	( 4'sd 4) * $signed(input_fmap_63[15:0]) +
	( 4'sd 5) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 4'sd 7) * $signed(input_fmap_67[15:0]) +
	( 3'sd 2) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_70[15:0]) +
	( 2'sd 1) * $signed(input_fmap_74[15:0]) +
	( 3'sd 2) * $signed(input_fmap_75[15:0]) +
	( 2'sd 1) * $signed(input_fmap_76[15:0]) +
	( 4'sd 7) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 3'sd 2) * $signed(input_fmap_80[15:0]) +
	( 4'sd 4) * $signed(input_fmap_81[15:0]) +
	( 4'sd 5) * $signed(input_fmap_82[15:0]) +
	( 4'sd 5) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 3'sd 3) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 3'sd 2) * $signed(input_fmap_88[15:0]) +
	( 2'sd 1) * $signed(input_fmap_89[15:0]) +
	( 4'sd 4) * $signed(input_fmap_90[15:0]) +
	( 4'sd 4) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 4'sd 4) * $signed(input_fmap_93[15:0]) +
	( 4'sd 4) * $signed(input_fmap_94[15:0]) +
	( 4'sd 7) * $signed(input_fmap_95[15:0]) +
	( 4'sd 7) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 6) * $signed(input_fmap_98[15:0]) +
	( 5'sd 8) * $signed(input_fmap_99[15:0]) +
	( 4'sd 4) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 4'sd 6) * $signed(input_fmap_102[15:0]) +
	( 4'sd 4) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 6) * $signed(input_fmap_105[15:0]) +
	( 2'sd 1) * $signed(input_fmap_106[15:0]) +
	( 3'sd 2) * $signed(input_fmap_107[15:0]) +
	( 4'sd 7) * $signed(input_fmap_108[15:0]) +
	( 4'sd 6) * $signed(input_fmap_109[15:0]) +
	( 4'sd 6) * $signed(input_fmap_111[15:0]) +
	( 4'sd 6) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 2'sd 1) * $signed(input_fmap_115[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 2'sd 1) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_119[15:0]) +
	( 2'sd 1) * $signed(input_fmap_120[15:0]) +
	( 4'sd 5) * $signed(input_fmap_121[15:0]) +
	( 4'sd 4) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_123[15:0]) +
	( 3'sd 3) * $signed(input_fmap_124[15:0]) +
	( 2'sd 1) * $signed(input_fmap_125[15:0]) +
	( 4'sd 5) * $signed(input_fmap_126[15:0]) +
	( 3'sd 2) * $signed(input_fmap_127[15:0]) +
	( 3'sd 3) * $signed(input_fmap_128[15:0]) +
	( 2'sd 1) * $signed(input_fmap_129[15:0]) +
	( 4'sd 4) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 4'sd 4) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 5'sd 8) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 3'sd 2) * $signed(input_fmap_136[15:0]) +
	( 4'sd 7) * $signed(input_fmap_137[15:0]) +
	( 3'sd 3) * $signed(input_fmap_138[15:0]) +
	( 2'sd 1) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 4'sd 4) * $signed(input_fmap_141[15:0]) +
	( 4'sd 6) * $signed(input_fmap_142[15:0]) +
	( 3'sd 2) * $signed(input_fmap_143[15:0]) +
	( 3'sd 3) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 4'sd 7) * $signed(input_fmap_146[15:0]) +
	( 3'sd 3) * $signed(input_fmap_147[15:0]) +
	( 4'sd 4) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 4'sd 4) * $signed(input_fmap_150[15:0]) +
	( 4'sd 4) * $signed(input_fmap_151[15:0]) +
	( 3'sd 2) * $signed(input_fmap_152[15:0]) +
	( 4'sd 7) * $signed(input_fmap_153[15:0]) +
	( 3'sd 2) * $signed(input_fmap_154[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 4) * $signed(input_fmap_157[15:0]) +
	( 2'sd 1) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 5'sd 8) * $signed(input_fmap_160[15:0]) +
	( 3'sd 2) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 3'sd 2) * $signed(input_fmap_163[15:0]) +
	( 3'sd 3) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 4'sd 4) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 3'sd 2) * $signed(input_fmap_168[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_170[15:0]) +
	( 4'sd 6) * $signed(input_fmap_171[15:0]) +
	( 4'sd 4) * $signed(input_fmap_172[15:0]) +
	( 3'sd 3) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 3'sd 2) * $signed(input_fmap_175[15:0]) +
	( 4'sd 7) * $signed(input_fmap_176[15:0]) +
	( 4'sd 7) * $signed(input_fmap_177[15:0]) +
	( 4'sd 6) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_182[15:0]) +
	( 2'sd 1) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 2'sd 1) * $signed(input_fmap_186[15:0]) +
	( 3'sd 3) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 3'sd 2) * $signed(input_fmap_189[15:0]) +
	( 4'sd 4) * $signed(input_fmap_190[15:0]) +
	( 5'sd 8) * $signed(input_fmap_191[15:0]) +
	( 4'sd 4) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 5) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 3'sd 3) * $signed(input_fmap_198[15:0]) +
	( 4'sd 4) * $signed(input_fmap_199[15:0]) +
	( 4'sd 7) * $signed(input_fmap_200[15:0]) +
	( 4'sd 6) * $signed(input_fmap_201[15:0]) +
	( 2'sd 1) * $signed(input_fmap_202[15:0]) +
	( 4'sd 6) * $signed(input_fmap_203[15:0]) +
	( 4'sd 7) * $signed(input_fmap_204[15:0]) +
	( 4'sd 7) * $signed(input_fmap_205[15:0]) +
	( 4'sd 5) * $signed(input_fmap_206[15:0]) +
	( 3'sd 3) * $signed(input_fmap_208[15:0]) +
	( 4'sd 6) * $signed(input_fmap_210[15:0]) +
	( 5'sd 8) * $signed(input_fmap_211[15:0]) +
	( 4'sd 4) * $signed(input_fmap_212[15:0]) +
	( 3'sd 2) * $signed(input_fmap_213[15:0]) +
	( 3'sd 2) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 4) * $signed(input_fmap_219[15:0]) +
	( 3'sd 2) * $signed(input_fmap_220[15:0]) +
	( 4'sd 5) * $signed(input_fmap_221[15:0]) +
	( 3'sd 2) * $signed(input_fmap_223[15:0]) +
	( 4'sd 4) * $signed(input_fmap_224[15:0]) +
	( 4'sd 6) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_227[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 3'sd 2) * $signed(input_fmap_230[15:0]) +
	( 4'sd 6) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 4'sd 5) * $signed(input_fmap_233[15:0]) +
	( 4'sd 4) * $signed(input_fmap_234[15:0]) +
	( 3'sd 3) * $signed(input_fmap_236[15:0]) +
	( 4'sd 7) * $signed(input_fmap_237[15:0]) +
	( 4'sd 6) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 3'sd 2) * $signed(input_fmap_240[15:0]) +
	( 3'sd 2) * $signed(input_fmap_241[15:0]) +
	( 4'sd 6) * $signed(input_fmap_242[15:0]) +
	( 2'sd 1) * $signed(input_fmap_243[15:0]) +
	( 4'sd 6) * $signed(input_fmap_244[15:0]) +
	( 4'sd 7) * $signed(input_fmap_245[15:0]) +
	( 4'sd 6) * $signed(input_fmap_246[15:0]) +
	( 3'sd 3) * $signed(input_fmap_247[15:0]) +
	( 3'sd 2) * $signed(input_fmap_248[15:0]) +
	( 5'sd 8) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 5) * $signed(input_fmap_254[15:0]) +
	( 4'sd 7) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_254;
assign conv_mac_254 = 
	( 5'sd 8) * $signed(input_fmap_0[15:0]) +
	( 5'sd 8) * $signed(input_fmap_1[15:0]) +
	( 4'sd 5) * $signed(input_fmap_2[15:0]) +
	( 4'sd 6) * $signed(input_fmap_3[15:0]) +
	( 5'sd 8) * $signed(input_fmap_4[15:0]) +
	( 3'sd 3) * $signed(input_fmap_5[15:0]) +
	( 4'sd 6) * $signed(input_fmap_6[15:0]) +
	( 4'sd 6) * $signed(input_fmap_7[15:0]) +
	( 3'sd 2) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 2'sd 1) * $signed(input_fmap_10[15:0]) +
	( 4'sd 6) * $signed(input_fmap_11[15:0]) +
	( 3'sd 3) * $signed(input_fmap_12[15:0]) +
	( 3'sd 3) * $signed(input_fmap_13[15:0]) +
	( 4'sd 7) * $signed(input_fmap_14[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 2'sd 1) * $signed(input_fmap_18[15:0]) +
	( 3'sd 3) * $signed(input_fmap_19[15:0]) +
	( 4'sd 6) * $signed(input_fmap_20[15:0]) +
	( 3'sd 3) * $signed(input_fmap_21[15:0]) +
	( 4'sd 4) * $signed(input_fmap_22[15:0]) +
	( 2'sd 1) * $signed(input_fmap_23[15:0]) +
	( 4'sd 7) * $signed(input_fmap_24[15:0]) +
	( 4'sd 5) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 6) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 4'sd 6) * $signed(input_fmap_30[15:0]) +
	( 2'sd 1) * $signed(input_fmap_31[15:0]) +
	( 3'sd 3) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 4'sd 6) * $signed(input_fmap_38[15:0]) +
	( 4'sd 7) * $signed(input_fmap_39[15:0]) +
	( 4'sd 6) * $signed(input_fmap_40[15:0]) +
	( 2'sd 1) * $signed(input_fmap_42[15:0]) +
	( 3'sd 2) * $signed(input_fmap_43[15:0]) +
	( 3'sd 2) * $signed(input_fmap_44[15:0]) +
	( 4'sd 4) * $signed(input_fmap_45[15:0]) +
	( 4'sd 5) * $signed(input_fmap_46[15:0]) +
	( 4'sd 5) * $signed(input_fmap_47[15:0]) +
	( 4'sd 6) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_49[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 2'sd 1) * $signed(input_fmap_51[15:0]) +
	( 4'sd 5) * $signed(input_fmap_52[15:0]) +
	( 4'sd 4) * $signed(input_fmap_53[15:0]) +
	( 4'sd 7) * $signed(input_fmap_54[15:0]) +
	( 3'sd 3) * $signed(input_fmap_55[15:0]) +
	( 3'sd 3) * $signed(input_fmap_56[15:0]) +
	( 2'sd 1) * $signed(input_fmap_57[15:0]) +
	( 2'sd 1) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 4'sd 6) * $signed(input_fmap_61[15:0]) +
	( 5'sd 8) * $signed(input_fmap_62[15:0]) +
	( 4'sd 5) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 4'sd 4) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 3'sd 3) * $signed(input_fmap_68[15:0]) +
	( 4'sd 7) * $signed(input_fmap_69[15:0]) +
	( 4'sd 6) * $signed(input_fmap_70[15:0]) +
	( 3'sd 2) * $signed(input_fmap_71[15:0]) +
	( 5'sd 8) * $signed(input_fmap_72[15:0]) +
	( 4'sd 7) * $signed(input_fmap_73[15:0]) +
	( 3'sd 3) * $signed(input_fmap_74[15:0]) +
	( 2'sd 1) * $signed(input_fmap_75[15:0]) +
	( 4'sd 7) * $signed(input_fmap_76[15:0]) +
	( 3'sd 3) * $signed(input_fmap_77[15:0]) +
	( 3'sd 2) * $signed(input_fmap_78[15:0]) +
	( 4'sd 7) * $signed(input_fmap_79[15:0]) +
	( 4'sd 5) * $signed(input_fmap_80[15:0]) +
	( 2'sd 1) * $signed(input_fmap_81[15:0]) +
	( 5'sd 8) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 2'sd 1) * $signed(input_fmap_84[15:0]) +
	( 3'sd 2) * $signed(input_fmap_85[15:0]) +
	( 2'sd 1) * $signed(input_fmap_86[15:0]) +
	( 5'sd 8) * $signed(input_fmap_87[15:0]) +
	( 4'sd 7) * $signed(input_fmap_88[15:0]) +
	( 5'sd 8) * $signed(input_fmap_89[15:0]) +
	( 3'sd 2) * $signed(input_fmap_90[15:0]) +
	( 4'sd 6) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 3'sd 3) * $signed(input_fmap_93[15:0]) +
	( 3'sd 2) * $signed(input_fmap_94[15:0]) +
	( 2'sd 1) * $signed(input_fmap_95[15:0]) +
	( 4'sd 6) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 3'sd 2) * $signed(input_fmap_98[15:0]) +
	( 3'sd 2) * $signed(input_fmap_99[15:0]) +
	( 5'sd 8) * $signed(input_fmap_100[15:0]) +
	( 4'sd 6) * $signed(input_fmap_101[15:0]) +
	( 2'sd 1) * $signed(input_fmap_102[15:0]) +
	( 3'sd 3) * $signed(input_fmap_103[15:0]) +
	( 4'sd 4) * $signed(input_fmap_104[15:0]) +
	( 3'sd 2) * $signed(input_fmap_105[15:0]) +
	( 3'sd 3) * $signed(input_fmap_106[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 3'sd 2) * $signed(input_fmap_108[15:0]) +
	( 4'sd 4) * $signed(input_fmap_109[15:0]) +
	( 3'sd 3) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 4) * $signed(input_fmap_113[15:0]) +
	( 4'sd 4) * $signed(input_fmap_114[15:0]) +
	( 4'sd 4) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 5) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 2) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 4'sd 5) * $signed(input_fmap_122[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 7) * $signed(input_fmap_125[15:0]) +
	( 4'sd 7) * $signed(input_fmap_126[15:0]) +
	( 3'sd 3) * $signed(input_fmap_127[15:0]) +
	( 4'sd 7) * $signed(input_fmap_128[15:0]) +
	( 4'sd 4) * $signed(input_fmap_129[15:0]) +
	( 3'sd 3) * $signed(input_fmap_130[15:0]) +
	( 5'sd 8) * $signed(input_fmap_131[15:0]) +
	( 4'sd 5) * $signed(input_fmap_132[15:0]) +
	( 3'sd 2) * $signed(input_fmap_133[15:0]) +
	( 3'sd 3) * $signed(input_fmap_134[15:0]) +
	( 5'sd 8) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_136[15:0]) +
	( 3'sd 3) * $signed(input_fmap_137[15:0]) +
	( 2'sd 1) * $signed(input_fmap_138[15:0]) +
	( 4'sd 4) * $signed(input_fmap_139[15:0]) +
	( 4'sd 6) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_143[15:0]) +
	( 3'sd 2) * $signed(input_fmap_144[15:0]) +
	( 4'sd 6) * $signed(input_fmap_145[15:0]) +
	( 2'sd 1) * $signed(input_fmap_146[15:0]) +
	( 4'sd 7) * $signed(input_fmap_147[15:0]) +
	( 5'sd 8) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 2'sd 1) * $signed(input_fmap_152[15:0]) +
	( 3'sd 2) * $signed(input_fmap_153[15:0]) +
	( 4'sd 7) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 3'sd 2) * $signed(input_fmap_156[15:0]) +
	( 5'sd 8) * $signed(input_fmap_157[15:0]) +
	( 3'sd 3) * $signed(input_fmap_158[15:0]) +
	( 5'sd 8) * $signed(input_fmap_159[15:0]) +
	( 4'sd 6) * $signed(input_fmap_160[15:0]) +
	( 4'sd 6) * $signed(input_fmap_161[15:0]) +
	( 4'sd 6) * $signed(input_fmap_162[15:0]) +
	( 4'sd 5) * $signed(input_fmap_163[15:0]) +
	( 3'sd 2) * $signed(input_fmap_164[15:0]) +
	( 4'sd 7) * $signed(input_fmap_165[15:0]) +
	( 4'sd 5) * $signed(input_fmap_166[15:0]) +
	( 3'sd 3) * $signed(input_fmap_167[15:0]) +
	( 4'sd 7) * $signed(input_fmap_169[15:0]) +
	( 4'sd 7) * $signed(input_fmap_170[15:0]) +
	( 5'sd 8) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 7) * $signed(input_fmap_173[15:0]) +
	( 4'sd 4) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 2'sd 1) * $signed(input_fmap_176[15:0]) +
	( 2'sd 1) * $signed(input_fmap_177[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 2'sd 1) * $signed(input_fmap_179[15:0]) +
	( 5'sd 8) * $signed(input_fmap_180[15:0]) +
	( 4'sd 5) * $signed(input_fmap_181[15:0]) +
	( 4'sd 7) * $signed(input_fmap_182[15:0]) +
	( 4'sd 7) * $signed(input_fmap_183[15:0]) +
	( 4'sd 6) * $signed(input_fmap_184[15:0]) +
	( 2'sd 1) * $signed(input_fmap_185[15:0]) +
	( 3'sd 3) * $signed(input_fmap_186[15:0]) +
	( 4'sd 4) * $signed(input_fmap_187[15:0]) +
	( 4'sd 6) * $signed(input_fmap_188[15:0]) +
	( 4'sd 4) * $signed(input_fmap_189[15:0]) +
	( 5'sd 8) * $signed(input_fmap_190[15:0]) +
	( 4'sd 5) * $signed(input_fmap_191[15:0]) +
	( 5'sd 8) * $signed(input_fmap_192[15:0]) +
	( 4'sd 5) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 7) * $signed(input_fmap_195[15:0]) +
	( 4'sd 5) * $signed(input_fmap_196[15:0]) +
	( 4'sd 7) * $signed(input_fmap_197[15:0]) +
	( 2'sd 1) * $signed(input_fmap_198[15:0]) +
	( 4'sd 5) * $signed(input_fmap_199[15:0]) +
	( 4'sd 5) * $signed(input_fmap_200[15:0]) +
	( 4'sd 4) * $signed(input_fmap_201[15:0]) +
	( 4'sd 6) * $signed(input_fmap_202[15:0]) +
	( 2'sd 1) * $signed(input_fmap_203[15:0]) +
	( 3'sd 2) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 4) * $signed(input_fmap_206[15:0]) +
	( 3'sd 2) * $signed(input_fmap_207[15:0]) +
	( 4'sd 5) * $signed(input_fmap_208[15:0]) +
	( 3'sd 3) * $signed(input_fmap_209[15:0]) +
	( 3'sd 2) * $signed(input_fmap_210[15:0]) +
	( 4'sd 6) * $signed(input_fmap_211[15:0]) +
	( 3'sd 2) * $signed(input_fmap_212[15:0]) +
	( 4'sd 7) * $signed(input_fmap_213[15:0]) +
	( 4'sd 4) * $signed(input_fmap_214[15:0]) +
	( 4'sd 7) * $signed(input_fmap_215[15:0]) +
	( 3'sd 2) * $signed(input_fmap_216[15:0]) +
	( 4'sd 4) * $signed(input_fmap_217[15:0]) +
	( 4'sd 4) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 3'sd 3) * $signed(input_fmap_220[15:0]) +
	( 4'sd 6) * $signed(input_fmap_221[15:0]) +
	( 4'sd 4) * $signed(input_fmap_222[15:0]) +
	( 4'sd 7) * $signed(input_fmap_224[15:0]) +
	( 3'sd 2) * $signed(input_fmap_225[15:0]) +
	( 4'sd 6) * $signed(input_fmap_226[15:0]) +
	( 3'sd 3) * $signed(input_fmap_228[15:0]) +
	( 4'sd 5) * $signed(input_fmap_229[15:0]) +
	( 3'sd 3) * $signed(input_fmap_231[15:0]) +
	( 4'sd 7) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 4'sd 6) * $signed(input_fmap_234[15:0]) +
	( 4'sd 6) * $signed(input_fmap_235[15:0]) +
	( 4'sd 7) * $signed(input_fmap_236[15:0]) +
	( 4'sd 4) * $signed(input_fmap_237[15:0]) +
	( 3'sd 2) * $signed(input_fmap_239[15:0]) +
	( 2'sd 1) * $signed(input_fmap_241[15:0]) +
	( 4'sd 7) * $signed(input_fmap_242[15:0]) +
	( 4'sd 6) * $signed(input_fmap_243[15:0]) +
	( 4'sd 5) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 4'sd 4) * $signed(input_fmap_246[15:0]) +
	( 5'sd 8) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 3'sd 2) * $signed(input_fmap_250[15:0]) +
	( 2'sd 1) * $signed(input_fmap_251[15:0]) +
	( 5'sd 8) * $signed(input_fmap_252[15:0]) +
	( 3'sd 3) * $signed(input_fmap_253[15:0]) +
	( 4'sd 6) * $signed(input_fmap_254[15:0]) +
	( 3'sd 3) * $signed(input_fmap_255[15:0]);

logic signed [31:0] conv_mac_255;
assign conv_mac_255 = 
	( 3'sd 2) * $signed(input_fmap_0[15:0]) +
	( 4'sd 6) * $signed(input_fmap_1[15:0]) +
	( 3'sd 3) * $signed(input_fmap_2[15:0]) +
	( 3'sd 2) * $signed(input_fmap_3[15:0]) +
	( 2'sd 1) * $signed(input_fmap_4[15:0]) +
	( 4'sd 5) * $signed(input_fmap_6[15:0]) +
	( 4'sd 7) * $signed(input_fmap_7[15:0]) +
	( 3'sd 3) * $signed(input_fmap_8[15:0]) +
	( 3'sd 2) * $signed(input_fmap_9[15:0]) +
	( 3'sd 3) * $signed(input_fmap_10[15:0]) +
	( 3'sd 3) * $signed(input_fmap_11[15:0]) +
	( 4'sd 4) * $signed(input_fmap_12[15:0]) +
	( 3'sd 2) * $signed(input_fmap_14[15:0]) +
	( 2'sd 1) * $signed(input_fmap_15[15:0]) +
	( 4'sd 6) * $signed(input_fmap_16[15:0]) +
	( 4'sd 5) * $signed(input_fmap_17[15:0]) +
	( 5'sd 8) * $signed(input_fmap_18[15:0]) +
	( 2'sd 1) * $signed(input_fmap_19[15:0]) +
	( 5'sd 8) * $signed(input_fmap_20[15:0]) +
	( 2'sd 1) * $signed(input_fmap_21[15:0]) +
	( 3'sd 2) * $signed(input_fmap_22[15:0]) +
	( 4'sd 5) * $signed(input_fmap_23[15:0]) +
	( 4'sd 4) * $signed(input_fmap_24[15:0]) +
	( 3'sd 3) * $signed(input_fmap_25[15:0]) +
	( 4'sd 5) * $signed(input_fmap_26[15:0]) +
	( 3'sd 2) * $signed(input_fmap_27[15:0]) +
	( 4'sd 4) * $signed(input_fmap_28[15:0]) +
	( 4'sd 5) * $signed(input_fmap_29[15:0]) +
	( 2'sd 1) * $signed(input_fmap_30[15:0]) +
	( 4'sd 4) * $signed(input_fmap_31[15:0]) +
	( 4'sd 4) * $signed(input_fmap_32[15:0]) +
	( 2'sd 1) * $signed(input_fmap_33[15:0]) +
	( 2'sd 1) * $signed(input_fmap_34[15:0]) +
	( 4'sd 5) * $signed(input_fmap_35[15:0]) +
	( 2'sd 1) * $signed(input_fmap_36[15:0]) +
	( 4'sd 6) * $signed(input_fmap_37[15:0]) +
	( 3'sd 3) * $signed(input_fmap_38[15:0]) +
	( 3'sd 2) * $signed(input_fmap_39[15:0]) +
	( 3'sd 2) * $signed(input_fmap_40[15:0]) +
	( 4'sd 6) * $signed(input_fmap_41[15:0]) +
	( 4'sd 4) * $signed(input_fmap_42[15:0]) +
	( 4'sd 7) * $signed(input_fmap_43[15:0]) +
	( 4'sd 4) * $signed(input_fmap_44[15:0]) +
	( 4'sd 7) * $signed(input_fmap_45[15:0]) +
	( 3'sd 2) * $signed(input_fmap_46[15:0]) +
	( 3'sd 2) * $signed(input_fmap_47[15:0]) +
	( 3'sd 2) * $signed(input_fmap_48[15:0]) +
	( 3'sd 2) * $signed(input_fmap_50[15:0]) +
	( 4'sd 6) * $signed(input_fmap_51[15:0]) +
	( 2'sd 1) * $signed(input_fmap_53[15:0]) +
	( 4'sd 4) * $signed(input_fmap_54[15:0]) +
	( 2'sd 1) * $signed(input_fmap_55[15:0]) +
	( 4'sd 5) * $signed(input_fmap_56[15:0]) +
	( 3'sd 3) * $signed(input_fmap_57[15:0]) +
	( 4'sd 4) * $signed(input_fmap_58[15:0]) +
	( 4'sd 5) * $signed(input_fmap_59[15:0]) +
	( 2'sd 1) * $signed(input_fmap_60[15:0]) +
	( 2'sd 1) * $signed(input_fmap_61[15:0]) +
	( 4'sd 4) * $signed(input_fmap_62[15:0]) +
	( 4'sd 6) * $signed(input_fmap_63[15:0]) +
	( 4'sd 4) * $signed(input_fmap_64[15:0]) +
	( 2'sd 1) * $signed(input_fmap_65[15:0]) +
	( 4'sd 7) * $signed(input_fmap_66[15:0]) +
	( 3'sd 3) * $signed(input_fmap_67[15:0]) +
	( 2'sd 1) * $signed(input_fmap_68[15:0]) +
	( 4'sd 4) * $signed(input_fmap_69[15:0]) +
	( 4'sd 5) * $signed(input_fmap_70[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 3'sd 3) * $signed(input_fmap_73[15:0]) +
	( 3'sd 2) * $signed(input_fmap_74[15:0]) +
	( 5'sd 8) * $signed(input_fmap_75[15:0]) +
	( 3'sd 2) * $signed(input_fmap_76[15:0]) +
	( 4'sd 4) * $signed(input_fmap_77[15:0]) +
	( 4'sd 7) * $signed(input_fmap_78[15:0]) +
	( 3'sd 3) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 3'sd 3) * $signed(input_fmap_81[15:0]) +
	( 4'sd 7) * $signed(input_fmap_82[15:0]) +
	( 3'sd 2) * $signed(input_fmap_83[15:0]) +
	( 4'sd 4) * $signed(input_fmap_84[15:0]) +
	( 4'sd 5) * $signed(input_fmap_85[15:0]) +
	( 4'sd 5) * $signed(input_fmap_86[15:0]) +
	( 4'sd 4) * $signed(input_fmap_87[15:0]) +
	( 2'sd 1) * $signed(input_fmap_88[15:0]) +
	( 4'sd 7) * $signed(input_fmap_89[15:0]) +
	( 2'sd 1) * $signed(input_fmap_90[15:0]) +
	( 4'sd 7) * $signed(input_fmap_91[15:0]) +
	( 2'sd 1) * $signed(input_fmap_92[15:0]) +
	( 2'sd 1) * $signed(input_fmap_93[15:0]) +
	( 4'sd 7) * $signed(input_fmap_94[15:0]) +
	( 4'sd 6) * $signed(input_fmap_95[15:0]) +
	( 3'sd 3) * $signed(input_fmap_96[15:0]) +
	( 3'sd 3) * $signed(input_fmap_97[15:0]) +
	( 4'sd 4) * $signed(input_fmap_98[15:0]) +
	( 4'sd 7) * $signed(input_fmap_99[15:0]) +
	( 3'sd 3) * $signed(input_fmap_100[15:0]) +
	( 4'sd 4) * $signed(input_fmap_101[15:0]) +
	( 4'sd 5) * $signed(input_fmap_102[15:0]) +
	( 4'sd 5) * $signed(input_fmap_103[15:0]) +
	( 4'sd 7) * $signed(input_fmap_104[15:0]) +
	( 4'sd 4) * $signed(input_fmap_105[15:0]) +
	( 4'sd 6) * $signed(input_fmap_107[15:0]) +
	( 2'sd 1) * $signed(input_fmap_108[15:0]) +
	( 3'sd 2) * $signed(input_fmap_109[15:0]) +
	( 3'sd 2) * $signed(input_fmap_110[15:0]) +
	( 4'sd 4) * $signed(input_fmap_111[15:0]) +
	( 4'sd 7) * $signed(input_fmap_112[15:0]) +
	( 2'sd 1) * $signed(input_fmap_113[15:0]) +
	( 4'sd 6) * $signed(input_fmap_114[15:0]) +
	( 4'sd 7) * $signed(input_fmap_116[15:0]) +
	( 4'sd 5) * $signed(input_fmap_117[15:0]) +
	( 4'sd 7) * $signed(input_fmap_118[15:0]) +
	( 4'sd 4) * $signed(input_fmap_119[15:0]) +
	( 3'sd 3) * $signed(input_fmap_120[15:0]) +
	( 4'sd 4) * $signed(input_fmap_121[15:0]) +
	( 3'sd 3) * $signed(input_fmap_122[15:0]) +
	( 4'sd 5) * $signed(input_fmap_123[15:0]) +
	( 4'sd 7) * $signed(input_fmap_124[15:0]) +
	( 4'sd 6) * $signed(input_fmap_125[15:0]) +
	( 4'sd 4) * $signed(input_fmap_126[15:0]) +
	( 2'sd 1) * $signed(input_fmap_127[15:0]) +
	( 4'sd 4) * $signed(input_fmap_128[15:0]) +
	( 5'sd 8) * $signed(input_fmap_129[15:0]) +
	( 4'sd 7) * $signed(input_fmap_130[15:0]) +
	( 4'sd 4) * $signed(input_fmap_131[15:0]) +
	( 2'sd 1) * $signed(input_fmap_132[15:0]) +
	( 4'sd 6) * $signed(input_fmap_133[15:0]) +
	( 4'sd 4) * $signed(input_fmap_134[15:0]) +
	( 4'sd 4) * $signed(input_fmap_135[15:0]) +
	( 4'sd 5) * $signed(input_fmap_137[15:0]) +
	( 5'sd 8) * $signed(input_fmap_138[15:0]) +
	( 4'sd 5) * $signed(input_fmap_139[15:0]) +
	( 3'sd 2) * $signed(input_fmap_140[15:0]) +
	( 2'sd 1) * $signed(input_fmap_141[15:0]) +
	( 4'sd 5) * $signed(input_fmap_142[15:0]) +
	( 4'sd 7) * $signed(input_fmap_143[15:0]) +
	( 2'sd 1) * $signed(input_fmap_144[15:0]) +
	( 4'sd 7) * $signed(input_fmap_145[15:0]) +
	( 3'sd 2) * $signed(input_fmap_146[15:0]) +
	( 4'sd 4) * $signed(input_fmap_147[15:0]) +
	( 3'sd 2) * $signed(input_fmap_148[15:0]) +
	( 4'sd 6) * $signed(input_fmap_149[15:0]) +
	( 3'sd 2) * $signed(input_fmap_150[15:0]) +
	( 4'sd 6) * $signed(input_fmap_151[15:0]) +
	( 5'sd 8) * $signed(input_fmap_152[15:0]) +
	( 5'sd 8) * $signed(input_fmap_153[15:0]) +
	( 5'sd 8) * $signed(input_fmap_154[15:0]) +
	( 3'sd 3) * $signed(input_fmap_155[15:0]) +
	( 4'sd 5) * $signed(input_fmap_156[15:0]) +
	( 4'sd 7) * $signed(input_fmap_157[15:0]) +
	( 4'sd 6) * $signed(input_fmap_158[15:0]) +
	( 3'sd 2) * $signed(input_fmap_159[15:0]) +
	( 4'sd 7) * $signed(input_fmap_160[15:0]) +
	( 4'sd 4) * $signed(input_fmap_161[15:0]) +
	( 4'sd 5) * $signed(input_fmap_162[15:0]) +
	( 4'sd 7) * $signed(input_fmap_163[15:0]) +
	( 2'sd 1) * $signed(input_fmap_164[15:0]) +
	( 2'sd 1) * $signed(input_fmap_165[15:0]) +
	( 5'sd 8) * $signed(input_fmap_166[15:0]) +
	( 4'sd 4) * $signed(input_fmap_167[15:0]) +
	( 5'sd 8) * $signed(input_fmap_168[15:0]) +
	( 5'sd 8) * $signed(input_fmap_169[15:0]) +
	( 4'sd 4) * $signed(input_fmap_171[15:0]) +
	( 4'sd 5) * $signed(input_fmap_172[15:0]) +
	( 4'sd 6) * $signed(input_fmap_173[15:0]) +
	( 2'sd 1) * $signed(input_fmap_174[15:0]) +
	( 4'sd 5) * $signed(input_fmap_175[15:0]) +
	( 5'sd 8) * $signed(input_fmap_176[15:0]) +
	( 3'sd 3) * $signed(input_fmap_178[15:0]) +
	( 4'sd 4) * $signed(input_fmap_179[15:0]) +
	( 3'sd 2) * $signed(input_fmap_180[15:0]) +
	( 4'sd 4) * $signed(input_fmap_181[15:0]) +
	( 4'sd 5) * $signed(input_fmap_182[15:0]) +
	( 4'sd 4) * $signed(input_fmap_183[15:0]) +
	( 2'sd 1) * $signed(input_fmap_184[15:0]) +
	( 4'sd 7) * $signed(input_fmap_185[15:0]) +
	( 4'sd 6) * $signed(input_fmap_186[15:0]) +
	( 2'sd 1) * $signed(input_fmap_187[15:0]) +
	( 4'sd 4) * $signed(input_fmap_188[15:0]) +
	( 4'sd 7) * $signed(input_fmap_189[15:0]) +
	( 2'sd 1) * $signed(input_fmap_190[15:0]) +
	( 2'sd 1) * $signed(input_fmap_191[15:0]) +
	( 4'sd 5) * $signed(input_fmap_192[15:0]) +
	( 4'sd 7) * $signed(input_fmap_193[15:0]) +
	( 2'sd 1) * $signed(input_fmap_194[15:0]) +
	( 4'sd 4) * $signed(input_fmap_195[15:0]) +
	( 3'sd 3) * $signed(input_fmap_196[15:0]) +
	( 4'sd 5) * $signed(input_fmap_197[15:0]) +
	( 3'sd 2) * $signed(input_fmap_198[15:0]) +
	( 4'sd 6) * $signed(input_fmap_199[15:0]) +
	( 3'sd 3) * $signed(input_fmap_200[15:0]) +
	( 2'sd 1) * $signed(input_fmap_201[15:0]) +
	( 3'sd 2) * $signed(input_fmap_202[15:0]) +
	( 4'sd 5) * $signed(input_fmap_203[15:0]) +
	( 4'sd 4) * $signed(input_fmap_204[15:0]) +
	( 4'sd 5) * $signed(input_fmap_205[15:0]) +
	( 4'sd 7) * $signed(input_fmap_206[15:0]) +
	( 4'sd 5) * $signed(input_fmap_207[15:0]) +
	( 5'sd 8) * $signed(input_fmap_208[15:0]) +
	( 2'sd 1) * $signed(input_fmap_209[15:0]) +
	( 4'sd 5) * $signed(input_fmap_210[15:0]) +
	( 4'sd 7) * $signed(input_fmap_211[15:0]) +
	( 3'sd 3) * $signed(input_fmap_212[15:0]) +
	( 5'sd 8) * $signed(input_fmap_214[15:0]) +
	( 3'sd 2) * $signed(input_fmap_215[15:0]) +
	( 2'sd 1) * $signed(input_fmap_216[15:0]) +
	( 3'sd 2) * $signed(input_fmap_217[15:0]) +
	( 2'sd 1) * $signed(input_fmap_218[15:0]) +
	( 4'sd 5) * $signed(input_fmap_219[15:0]) +
	( 4'sd 4) * $signed(input_fmap_221[15:0]) +
	( 5'sd 8) * $signed(input_fmap_222[15:0]) +
	( 3'sd 3) * $signed(input_fmap_223[15:0]) +
	( 2'sd 1) * $signed(input_fmap_224[15:0]) +
	( 4'sd 4) * $signed(input_fmap_225[15:0]) +
	( 2'sd 1) * $signed(input_fmap_226[15:0]) +
	( 2'sd 1) * $signed(input_fmap_227[15:0]) +
	( 3'sd 2) * $signed(input_fmap_228[15:0]) +
	( 2'sd 1) * $signed(input_fmap_229[15:0]) +
	( 4'sd 5) * $signed(input_fmap_230[15:0]) +
	( 4'sd 4) * $signed(input_fmap_231[15:0]) +
	( 4'sd 5) * $signed(input_fmap_232[15:0]) +
	( 2'sd 1) * $signed(input_fmap_233[15:0]) +
	( 3'sd 3) * $signed(input_fmap_234[15:0]) +
	( 4'sd 7) * $signed(input_fmap_235[15:0]) +
	( 3'sd 2) * $signed(input_fmap_236[15:0]) +
	( 3'sd 3) * $signed(input_fmap_237[15:0]) +
	( 3'sd 3) * $signed(input_fmap_238[15:0]) +
	( 4'sd 6) * $signed(input_fmap_239[15:0]) +
	( 4'sd 4) * $signed(input_fmap_241[15:0]) +
	( 4'sd 4) * $signed(input_fmap_242[15:0]) +
	( 4'sd 5) * $signed(input_fmap_243[15:0]) +
	( 5'sd 8) * $signed(input_fmap_244[15:0]) +
	( 4'sd 6) * $signed(input_fmap_245[15:0]) +
	( 3'sd 2) * $signed(input_fmap_246[15:0]) +
	( 4'sd 4) * $signed(input_fmap_247[15:0]) +
	( 2'sd 1) * $signed(input_fmap_248[15:0]) +
	( 4'sd 7) * $signed(input_fmap_249[15:0]) +
	( 2'sd 1) * $signed(input_fmap_250[15:0]) +
	( 3'sd 2) * $signed(input_fmap_251[15:0]) +
	( 4'sd 6) * $signed(input_fmap_252[15:0]) +
	( 5'sd 8) * $signed(input_fmap_253[15:0]) +
	( 2'sd 1) * $signed(input_fmap_254[15:0]) +
	( 3'sd 2) * $signed(input_fmap_255[15:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 5'd8;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 3'd3;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 2'd1;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 3'd3;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 3'd2;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 2'd1;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 3'd2;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 4'd6;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 4'd7;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 4'd6;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 4'd4;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 4'd4;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 2'd1;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 3'd3;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 4'd7;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 4'd5;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 2'd1;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 4'd7;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 3'd2;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 4'd6;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 4'd4;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 4'd6;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 4'd6;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 3'd2;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 3'd3;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 3'd2;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 4'd7;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 5'd8;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 3'd3;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 2'd1;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 3'd3;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 2'd1;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 4'd6;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 3'd2;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 4'd7;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 4'd5;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 4'd4;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 3'd2;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 2'd1;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 2'd1;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 3'd3;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 2'd1;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 5'd8;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 4'd6;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 4'd6;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 4'd5;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 4'd5;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 5'd8;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 4'd7;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 2'd1;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 2'd1;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 4'd6;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 3'd3;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 4'd7;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 4'd4;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 4'd7;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 4'd7;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 4'd4;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 2'd1;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 4'd4;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 2'd1;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 3'd2;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 4'd5;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 3'd2;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 3'd3;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 3'd3;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 3'd3;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 4'd5;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 4'd5;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 4'd6;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 4'd7;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 5'd8;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 4'd5;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 4'd5;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 2'd1;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 3'd2;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 4'd5;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 3'd2;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 4'd6;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 3'd2;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 4'd4;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 3'd3;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 3'd2;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 3'd2;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 3'd2;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 2'd1;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 3'd3;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 5'd8;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 4'd5;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 4'd5;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 4'd5;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 3'd2;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 4'd5;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 4'd6;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 4'd4;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 3'd3;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 3'd3;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 4'd5;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 4'd7;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 4'd4;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 4'd6;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 2'd1;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 4'd7;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 4'd4;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 3'd2;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 4'd4;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 4'd4;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 5'd8;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 2'd1;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 2'd1;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 4'd6;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 4'd5;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 4'd5;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 4'd5;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 4'd4;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 4'd5;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 3'd2;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 4'd7;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 4'd6;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 4'd5;
logic [31:0] bias_add_128;
assign bias_add_128 = conv_mac_128 + 3'd3;
logic [31:0] bias_add_129;
assign bias_add_129 = conv_mac_129 + 3'd2;
logic [31:0] bias_add_130;
assign bias_add_130 = conv_mac_130 + 2'd1;
logic [31:0] bias_add_131;
assign bias_add_131 = conv_mac_131 + 3'd3;
logic [31:0] bias_add_132;
assign bias_add_132 = conv_mac_132 + 4'd7;
logic [31:0] bias_add_133;
assign bias_add_133 = conv_mac_133 + 4'd4;
logic [31:0] bias_add_134;
assign bias_add_134 = conv_mac_134 + 4'd4;
logic [31:0] bias_add_135;
assign bias_add_135 = conv_mac_135 + 4'd7;
logic [31:0] bias_add_136;
assign bias_add_136 = conv_mac_136 + 4'd7;
logic [31:0] bias_add_137;
assign bias_add_137 = conv_mac_137 + 5'd8;
logic [31:0] bias_add_138;
assign bias_add_138 = conv_mac_138 + 4'd5;
logic [31:0] bias_add_139;
assign bias_add_139 = conv_mac_139;
logic [31:0] bias_add_140;
assign bias_add_140 = conv_mac_140 + 3'd2;
logic [31:0] bias_add_141;
assign bias_add_141 = conv_mac_141 + 3'd2;
logic [31:0] bias_add_142;
assign bias_add_142 = conv_mac_142;
logic [31:0] bias_add_143;
assign bias_add_143 = conv_mac_143 + 5'd8;
logic [31:0] bias_add_144;
assign bias_add_144 = conv_mac_144 + 4'd4;
logic [31:0] bias_add_145;
assign bias_add_145 = conv_mac_145 + 3'd3;
logic [31:0] bias_add_146;
assign bias_add_146 = conv_mac_146 + 2'd1;
logic [31:0] bias_add_147;
assign bias_add_147 = conv_mac_147 + 4'd7;
logic [31:0] bias_add_148;
assign bias_add_148 = conv_mac_148 + 4'd5;
logic [31:0] bias_add_149;
assign bias_add_149 = conv_mac_149 + 4'd7;
logic [31:0] bias_add_150;
assign bias_add_150 = conv_mac_150 + 2'd1;
logic [31:0] bias_add_151;
assign bias_add_151 = conv_mac_151 + 4'd4;
logic [31:0] bias_add_152;
assign bias_add_152 = conv_mac_152 + 4'd4;
logic [31:0] bias_add_153;
assign bias_add_153 = conv_mac_153 + 4'd7;
logic [31:0] bias_add_154;
assign bias_add_154 = conv_mac_154 + 3'd3;
logic [31:0] bias_add_155;
assign bias_add_155 = conv_mac_155 + 3'd2;
logic [31:0] bias_add_156;
assign bias_add_156 = conv_mac_156 + 5'd8;
logic [31:0] bias_add_157;
assign bias_add_157 = conv_mac_157;
logic [31:0] bias_add_158;
assign bias_add_158 = conv_mac_158 + 3'd3;
logic [31:0] bias_add_159;
assign bias_add_159 = conv_mac_159 + 4'd5;
logic [31:0] bias_add_160;
assign bias_add_160 = conv_mac_160 + 4'd6;
logic [31:0] bias_add_161;
assign bias_add_161 = conv_mac_161 + 4'd4;
logic [31:0] bias_add_162;
assign bias_add_162 = conv_mac_162 + 4'd4;
logic [31:0] bias_add_163;
assign bias_add_163 = conv_mac_163 + 5'd8;
logic [31:0] bias_add_164;
assign bias_add_164 = conv_mac_164 + 4'd6;
logic [31:0] bias_add_165;
assign bias_add_165 = conv_mac_165 + 4'd7;
logic [31:0] bias_add_166;
assign bias_add_166 = conv_mac_166 + 2'd1;
logic [31:0] bias_add_167;
assign bias_add_167 = conv_mac_167 + 4'd6;
logic [31:0] bias_add_168;
assign bias_add_168 = conv_mac_168 + 4'd4;
logic [31:0] bias_add_169;
assign bias_add_169 = conv_mac_169 + 4'd6;
logic [31:0] bias_add_170;
assign bias_add_170 = conv_mac_170 + 4'd6;
logic [31:0] bias_add_171;
assign bias_add_171 = conv_mac_171 + 4'd5;
logic [31:0] bias_add_172;
assign bias_add_172 = conv_mac_172 + 4'd7;
logic [31:0] bias_add_173;
assign bias_add_173 = conv_mac_173 + 4'd6;
logic [31:0] bias_add_174;
assign bias_add_174 = conv_mac_174;
logic [31:0] bias_add_175;
assign bias_add_175 = conv_mac_175 + 4'd7;
logic [31:0] bias_add_176;
assign bias_add_176 = conv_mac_176 + 4'd6;
logic [31:0] bias_add_177;
assign bias_add_177 = conv_mac_177 + 2'd1;
logic [31:0] bias_add_178;
assign bias_add_178 = conv_mac_178 + 4'd6;
logic [31:0] bias_add_179;
assign bias_add_179 = conv_mac_179 + 4'd6;
logic [31:0] bias_add_180;
assign bias_add_180 = conv_mac_180 + 4'd6;
logic [31:0] bias_add_181;
assign bias_add_181 = conv_mac_181 + 4'd5;
logic [31:0] bias_add_182;
assign bias_add_182 = conv_mac_182 + 4'd4;
logic [31:0] bias_add_183;
assign bias_add_183 = conv_mac_183 + 5'd8;
logic [31:0] bias_add_184;
assign bias_add_184 = conv_mac_184 + 4'd4;
logic [31:0] bias_add_185;
assign bias_add_185 = conv_mac_185 + 4'd4;
logic [31:0] bias_add_186;
assign bias_add_186 = conv_mac_186 + 3'd3;
logic [31:0] bias_add_187;
assign bias_add_187 = conv_mac_187 + 4'd4;
logic [31:0] bias_add_188;
assign bias_add_188 = conv_mac_188 + 4'd7;
logic [31:0] bias_add_189;
assign bias_add_189 = conv_mac_189 + 3'd2;
logic [31:0] bias_add_190;
assign bias_add_190 = conv_mac_190;
logic [31:0] bias_add_191;
assign bias_add_191 = conv_mac_191;
logic [31:0] bias_add_192;
assign bias_add_192 = conv_mac_192 + 4'd5;
logic [31:0] bias_add_193;
assign bias_add_193 = conv_mac_193 + 4'd5;
logic [31:0] bias_add_194;
assign bias_add_194 = conv_mac_194 + 4'd5;
logic [31:0] bias_add_195;
assign bias_add_195 = conv_mac_195 + 2'd1;
logic [31:0] bias_add_196;
assign bias_add_196 = conv_mac_196 + 2'd1;
logic [31:0] bias_add_197;
assign bias_add_197 = conv_mac_197 + 5'd8;
logic [31:0] bias_add_198;
assign bias_add_198 = conv_mac_198 + 4'd4;
logic [31:0] bias_add_199;
assign bias_add_199 = conv_mac_199 + 3'd2;
logic [31:0] bias_add_200;
assign bias_add_200 = conv_mac_200 + 2'd1;
logic [31:0] bias_add_201;
assign bias_add_201 = conv_mac_201 + 2'd1;
logic [31:0] bias_add_202;
assign bias_add_202 = conv_mac_202 + 4'd6;
logic [31:0] bias_add_203;
assign bias_add_203 = conv_mac_203 + 2'd1;
logic [31:0] bias_add_204;
assign bias_add_204 = conv_mac_204 + 4'd7;
logic [31:0] bias_add_205;
assign bias_add_205 = conv_mac_205 + 4'd6;
logic [31:0] bias_add_206;
assign bias_add_206 = conv_mac_206 + 3'd3;
logic [31:0] bias_add_207;
assign bias_add_207 = conv_mac_207 + 3'd3;
logic [31:0] bias_add_208;
assign bias_add_208 = conv_mac_208 + 4'd7;
logic [31:0] bias_add_209;
assign bias_add_209 = conv_mac_209 + 4'd5;
logic [31:0] bias_add_210;
assign bias_add_210 = conv_mac_210 + 4'd6;
logic [31:0] bias_add_211;
assign bias_add_211 = conv_mac_211 + 4'd6;
logic [31:0] bias_add_212;
assign bias_add_212 = conv_mac_212;
logic [31:0] bias_add_213;
assign bias_add_213 = conv_mac_213 + 4'd5;
logic [31:0] bias_add_214;
assign bias_add_214 = conv_mac_214 + 4'd6;
logic [31:0] bias_add_215;
assign bias_add_215 = conv_mac_215 + 4'd5;
logic [31:0] bias_add_216;
assign bias_add_216 = conv_mac_216 + 4'd6;
logic [31:0] bias_add_217;
assign bias_add_217 = conv_mac_217 + 2'd1;
logic [31:0] bias_add_218;
assign bias_add_218 = conv_mac_218 + 5'd8;
logic [31:0] bias_add_219;
assign bias_add_219 = conv_mac_219 + 2'd1;
logic [31:0] bias_add_220;
assign bias_add_220 = conv_mac_220 + 2'd1;
logic [31:0] bias_add_221;
assign bias_add_221 = conv_mac_221 + 3'd2;
logic [31:0] bias_add_222;
assign bias_add_222 = conv_mac_222 + 4'd4;
logic [31:0] bias_add_223;
assign bias_add_223 = conv_mac_223 + 2'd1;
logic [31:0] bias_add_224;
assign bias_add_224 = conv_mac_224 + 4'd7;
logic [31:0] bias_add_225;
assign bias_add_225 = conv_mac_225 + 4'd6;
logic [31:0] bias_add_226;
assign bias_add_226 = conv_mac_226 + 3'd3;
logic [31:0] bias_add_227;
assign bias_add_227 = conv_mac_227 + 2'd1;
logic [31:0] bias_add_228;
assign bias_add_228 = conv_mac_228 + 3'd3;
logic [31:0] bias_add_229;
assign bias_add_229 = conv_mac_229 + 2'd1;
logic [31:0] bias_add_230;
assign bias_add_230 = conv_mac_230 + 3'd3;
logic [31:0] bias_add_231;
assign bias_add_231 = conv_mac_231 + 4'd7;
logic [31:0] bias_add_232;
assign bias_add_232 = conv_mac_232 + 3'd3;
logic [31:0] bias_add_233;
assign bias_add_233 = conv_mac_233 + 4'd6;
logic [31:0] bias_add_234;
assign bias_add_234 = conv_mac_234 + 2'd1;
logic [31:0] bias_add_235;
assign bias_add_235 = conv_mac_235 + 4'd7;
logic [31:0] bias_add_236;
assign bias_add_236 = conv_mac_236;
logic [31:0] bias_add_237;
assign bias_add_237 = conv_mac_237 + 5'd8;
logic [31:0] bias_add_238;
assign bias_add_238 = conv_mac_238 + 2'd1;
logic [31:0] bias_add_239;
assign bias_add_239 = conv_mac_239 + 4'd4;
logic [31:0] bias_add_240;
assign bias_add_240 = conv_mac_240 + 4'd6;
logic [31:0] bias_add_241;
assign bias_add_241 = conv_mac_241 + 2'd1;
logic [31:0] bias_add_242;
assign bias_add_242 = conv_mac_242 + 3'd3;
logic [31:0] bias_add_243;
assign bias_add_243 = conv_mac_243 + 2'd1;
logic [31:0] bias_add_244;
assign bias_add_244 = conv_mac_244 + 5'd8;
logic [31:0] bias_add_245;
assign bias_add_245 = conv_mac_245 + 4'd7;
logic [31:0] bias_add_246;
assign bias_add_246 = conv_mac_246 + 4'd4;
logic [31:0] bias_add_247;
assign bias_add_247 = conv_mac_247 + 5'd8;
logic [31:0] bias_add_248;
assign bias_add_248 = conv_mac_248 + 4'd4;
logic [31:0] bias_add_249;
assign bias_add_249 = conv_mac_249 + 4'd7;
logic [31:0] bias_add_250;
assign bias_add_250 = conv_mac_250 + 2'd1;
logic [31:0] bias_add_251;
assign bias_add_251 = conv_mac_251 + 4'd6;
logic [31:0] bias_add_252;
assign bias_add_252 = conv_mac_252 + 4'd6;
logic [31:0] bias_add_253;
assign bias_add_253 = conv_mac_253;
logic [31:0] bias_add_254;
assign bias_add_254 = conv_mac_254 + 3'd3;
logic [31:0] bias_add_255;
assign bias_add_255 = conv_mac_255 + 2'd1;

logic [15:0] relu_0;
assign relu_0[15:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[17:3]}} :'d6) : '0;
logic [15:0] relu_1;
assign relu_1[15:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[17:3]}} :'d6) : '0;
logic [15:0] relu_2;
assign relu_2[15:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[17:3]}} :'d6) : '0;
logic [15:0] relu_3;
assign relu_3[15:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[17:3]}} :'d6) : '0;
logic [15:0] relu_4;
assign relu_4[15:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[17:3]}} :'d6) : '0;
logic [15:0] relu_5;
assign relu_5[15:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[17:3]}} :'d6) : '0;
logic [15:0] relu_6;
assign relu_6[15:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[17:3]}} :'d6) : '0;
logic [15:0] relu_7;
assign relu_7[15:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[17:3]}} :'d6) : '0;
logic [15:0] relu_8;
assign relu_8[15:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[17:3]}} :'d6) : '0;
logic [15:0] relu_9;
assign relu_9[15:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[17:3]}} :'d6) : '0;
logic [15:0] relu_10;
assign relu_10[15:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[17:3]}} :'d6) : '0;
logic [15:0] relu_11;
assign relu_11[15:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[17:3]}} :'d6) : '0;
logic [15:0] relu_12;
assign relu_12[15:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[17:3]}} :'d6) : '0;
logic [15:0] relu_13;
assign relu_13[15:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[17:3]}} :'d6) : '0;
logic [15:0] relu_14;
assign relu_14[15:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[17:3]}} :'d6) : '0;
logic [15:0] relu_15;
assign relu_15[15:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[17:3]}} :'d6) : '0;
logic [15:0] relu_16;
assign relu_16[15:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[17:3]}} :'d6) : '0;
logic [15:0] relu_17;
assign relu_17[15:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[17:3]}} :'d6) : '0;
logic [15:0] relu_18;
assign relu_18[15:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[17:3]}} :'d6) : '0;
logic [15:0] relu_19;
assign relu_19[15:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[17:3]}} :'d6) : '0;
logic [15:0] relu_20;
assign relu_20[15:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[17:3]}} :'d6) : '0;
logic [15:0] relu_21;
assign relu_21[15:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[17:3]}} :'d6) : '0;
logic [15:0] relu_22;
assign relu_22[15:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[17:3]}} :'d6) : '0;
logic [15:0] relu_23;
assign relu_23[15:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[17:3]}} :'d6) : '0;
logic [15:0] relu_24;
assign relu_24[15:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[17:3]}} :'d6) : '0;
logic [15:0] relu_25;
assign relu_25[15:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[17:3]}} :'d6) : '0;
logic [15:0] relu_26;
assign relu_26[15:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[17:3]}} :'d6) : '0;
logic [15:0] relu_27;
assign relu_27[15:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[17:3]}} :'d6) : '0;
logic [15:0] relu_28;
assign relu_28[15:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[17:3]}} :'d6) : '0;
logic [15:0] relu_29;
assign relu_29[15:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[17:3]}} :'d6) : '0;
logic [15:0] relu_30;
assign relu_30[15:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[17:3]}} :'d6) : '0;
logic [15:0] relu_31;
assign relu_31[15:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[17:3]}} :'d6) : '0;
logic [15:0] relu_32;
assign relu_32[15:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[17:3]}} :'d6) : '0;
logic [15:0] relu_33;
assign relu_33[15:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[17:3]}} :'d6) : '0;
logic [15:0] relu_34;
assign relu_34[15:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[17:3]}} :'d6) : '0;
logic [15:0] relu_35;
assign relu_35[15:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[17:3]}} :'d6) : '0;
logic [15:0] relu_36;
assign relu_36[15:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[17:3]}} :'d6) : '0;
logic [15:0] relu_37;
assign relu_37[15:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[17:3]}} :'d6) : '0;
logic [15:0] relu_38;
assign relu_38[15:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[17:3]}} :'d6) : '0;
logic [15:0] relu_39;
assign relu_39[15:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[17:3]}} :'d6) : '0;
logic [15:0] relu_40;
assign relu_40[15:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[17:3]}} :'d6) : '0;
logic [15:0] relu_41;
assign relu_41[15:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[17:3]}} :'d6) : '0;
logic [15:0] relu_42;
assign relu_42[15:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[17:3]}} :'d6) : '0;
logic [15:0] relu_43;
assign relu_43[15:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[17:3]}} :'d6) : '0;
logic [15:0] relu_44;
assign relu_44[15:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[17:3]}} :'d6) : '0;
logic [15:0] relu_45;
assign relu_45[15:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[17:3]}} :'d6) : '0;
logic [15:0] relu_46;
assign relu_46[15:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[17:3]}} :'d6) : '0;
logic [15:0] relu_47;
assign relu_47[15:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[17:3]}} :'d6) : '0;
logic [15:0] relu_48;
assign relu_48[15:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[17:3]}} :'d6) : '0;
logic [15:0] relu_49;
assign relu_49[15:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[17:3]}} :'d6) : '0;
logic [15:0] relu_50;
assign relu_50[15:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[17:3]}} :'d6) : '0;
logic [15:0] relu_51;
assign relu_51[15:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[17:3]}} :'d6) : '0;
logic [15:0] relu_52;
assign relu_52[15:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[17:3]}} :'d6) : '0;
logic [15:0] relu_53;
assign relu_53[15:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[17:3]}} :'d6) : '0;
logic [15:0] relu_54;
assign relu_54[15:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[17:3]}} :'d6) : '0;
logic [15:0] relu_55;
assign relu_55[15:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[17:3]}} :'d6) : '0;
logic [15:0] relu_56;
assign relu_56[15:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[17:3]}} :'d6) : '0;
logic [15:0] relu_57;
assign relu_57[15:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[17:3]}} :'d6) : '0;
logic [15:0] relu_58;
assign relu_58[15:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[17:3]}} :'d6) : '0;
logic [15:0] relu_59;
assign relu_59[15:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[17:3]}} :'d6) : '0;
logic [15:0] relu_60;
assign relu_60[15:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[17:3]}} :'d6) : '0;
logic [15:0] relu_61;
assign relu_61[15:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[17:3]}} :'d6) : '0;
logic [15:0] relu_62;
assign relu_62[15:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[17:3]}} :'d6) : '0;
logic [15:0] relu_63;
assign relu_63[15:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[17:3]}} :'d6) : '0;
logic [15:0] relu_64;
assign relu_64[15:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[17:3]}} :'d6) : '0;
logic [15:0] relu_65;
assign relu_65[15:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[17:3]}} :'d6) : '0;
logic [15:0] relu_66;
assign relu_66[15:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[17:3]}} :'d6) : '0;
logic [15:0] relu_67;
assign relu_67[15:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[17:3]}} :'d6) : '0;
logic [15:0] relu_68;
assign relu_68[15:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[17:3]}} :'d6) : '0;
logic [15:0] relu_69;
assign relu_69[15:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[17:3]}} :'d6) : '0;
logic [15:0] relu_70;
assign relu_70[15:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[17:3]}} :'d6) : '0;
logic [15:0] relu_71;
assign relu_71[15:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[17:3]}} :'d6) : '0;
logic [15:0] relu_72;
assign relu_72[15:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[17:3]}} :'d6) : '0;
logic [15:0] relu_73;
assign relu_73[15:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[17:3]}} :'d6) : '0;
logic [15:0] relu_74;
assign relu_74[15:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[17:3]}} :'d6) : '0;
logic [15:0] relu_75;
assign relu_75[15:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[17:3]}} :'d6) : '0;
logic [15:0] relu_76;
assign relu_76[15:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[17:3]}} :'d6) : '0;
logic [15:0] relu_77;
assign relu_77[15:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[17:3]}} :'d6) : '0;
logic [15:0] relu_78;
assign relu_78[15:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[17:3]}} :'d6) : '0;
logic [15:0] relu_79;
assign relu_79[15:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[17:3]}} :'d6) : '0;
logic [15:0] relu_80;
assign relu_80[15:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[17:3]}} :'d6) : '0;
logic [15:0] relu_81;
assign relu_81[15:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[17:3]}} :'d6) : '0;
logic [15:0] relu_82;
assign relu_82[15:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[17:3]}} :'d6) : '0;
logic [15:0] relu_83;
assign relu_83[15:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[17:3]}} :'d6) : '0;
logic [15:0] relu_84;
assign relu_84[15:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[17:3]}} :'d6) : '0;
logic [15:0] relu_85;
assign relu_85[15:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[17:3]}} :'d6) : '0;
logic [15:0] relu_86;
assign relu_86[15:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[17:3]}} :'d6) : '0;
logic [15:0] relu_87;
assign relu_87[15:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[17:3]}} :'d6) : '0;
logic [15:0] relu_88;
assign relu_88[15:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[17:3]}} :'d6) : '0;
logic [15:0] relu_89;
assign relu_89[15:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[17:3]}} :'d6) : '0;
logic [15:0] relu_90;
assign relu_90[15:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[17:3]}} :'d6) : '0;
logic [15:0] relu_91;
assign relu_91[15:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[17:3]}} :'d6) : '0;
logic [15:0] relu_92;
assign relu_92[15:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[17:3]}} :'d6) : '0;
logic [15:0] relu_93;
assign relu_93[15:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[17:3]}} :'d6) : '0;
logic [15:0] relu_94;
assign relu_94[15:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[17:3]}} :'d6) : '0;
logic [15:0] relu_95;
assign relu_95[15:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[17:3]}} :'d6) : '0;
logic [15:0] relu_96;
assign relu_96[15:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[17:3]}} :'d6) : '0;
logic [15:0] relu_97;
assign relu_97[15:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[17:3]}} :'d6) : '0;
logic [15:0] relu_98;
assign relu_98[15:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[17:3]}} :'d6) : '0;
logic [15:0] relu_99;
assign relu_99[15:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[17:3]}} :'d6) : '0;
logic [15:0] relu_100;
assign relu_100[15:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[17:3]}} :'d6) : '0;
logic [15:0] relu_101;
assign relu_101[15:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[17:3]}} :'d6) : '0;
logic [15:0] relu_102;
assign relu_102[15:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[17:3]}} :'d6) : '0;
logic [15:0] relu_103;
assign relu_103[15:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[17:3]}} :'d6) : '0;
logic [15:0] relu_104;
assign relu_104[15:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[17:3]}} :'d6) : '0;
logic [15:0] relu_105;
assign relu_105[15:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[17:3]}} :'d6) : '0;
logic [15:0] relu_106;
assign relu_106[15:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[17:3]}} :'d6) : '0;
logic [15:0] relu_107;
assign relu_107[15:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[17:3]}} :'d6) : '0;
logic [15:0] relu_108;
assign relu_108[15:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[17:3]}} :'d6) : '0;
logic [15:0] relu_109;
assign relu_109[15:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[17:3]}} :'d6) : '0;
logic [15:0] relu_110;
assign relu_110[15:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[17:3]}} :'d6) : '0;
logic [15:0] relu_111;
assign relu_111[15:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[17:3]}} :'d6) : '0;
logic [15:0] relu_112;
assign relu_112[15:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[17:3]}} :'d6) : '0;
logic [15:0] relu_113;
assign relu_113[15:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[17:3]}} :'d6) : '0;
logic [15:0] relu_114;
assign relu_114[15:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[17:3]}} :'d6) : '0;
logic [15:0] relu_115;
assign relu_115[15:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[17:3]}} :'d6) : '0;
logic [15:0] relu_116;
assign relu_116[15:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[17:3]}} :'d6) : '0;
logic [15:0] relu_117;
assign relu_117[15:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[17:3]}} :'d6) : '0;
logic [15:0] relu_118;
assign relu_118[15:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[17:3]}} :'d6) : '0;
logic [15:0] relu_119;
assign relu_119[15:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[17:3]}} :'d6) : '0;
logic [15:0] relu_120;
assign relu_120[15:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[17:3]}} :'d6) : '0;
logic [15:0] relu_121;
assign relu_121[15:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[17:3]}} :'d6) : '0;
logic [15:0] relu_122;
assign relu_122[15:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[17:3]}} :'d6) : '0;
logic [15:0] relu_123;
assign relu_123[15:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[17:3]}} :'d6) : '0;
logic [15:0] relu_124;
assign relu_124[15:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[17:3]}} :'d6) : '0;
logic [15:0] relu_125;
assign relu_125[15:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[17:3]}} :'d6) : '0;
logic [15:0] relu_126;
assign relu_126[15:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[17:3]}} :'d6) : '0;
logic [15:0] relu_127;
assign relu_127[15:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[17:3]}} :'d6) : '0;
logic [15:0] relu_128;
assign relu_128[15:0] = (bias_add_128[31]==0) ? ((bias_add_128<3'd6) ? {{bias_add_128[31],bias_add_128[17:3]}} :'d6) : '0;
logic [15:0] relu_129;
assign relu_129[15:0] = (bias_add_129[31]==0) ? ((bias_add_129<3'd6) ? {{bias_add_129[31],bias_add_129[17:3]}} :'d6) : '0;
logic [15:0] relu_130;
assign relu_130[15:0] = (bias_add_130[31]==0) ? ((bias_add_130<3'd6) ? {{bias_add_130[31],bias_add_130[17:3]}} :'d6) : '0;
logic [15:0] relu_131;
assign relu_131[15:0] = (bias_add_131[31]==0) ? ((bias_add_131<3'd6) ? {{bias_add_131[31],bias_add_131[17:3]}} :'d6) : '0;
logic [15:0] relu_132;
assign relu_132[15:0] = (bias_add_132[31]==0) ? ((bias_add_132<3'd6) ? {{bias_add_132[31],bias_add_132[17:3]}} :'d6) : '0;
logic [15:0] relu_133;
assign relu_133[15:0] = (bias_add_133[31]==0) ? ((bias_add_133<3'd6) ? {{bias_add_133[31],bias_add_133[17:3]}} :'d6) : '0;
logic [15:0] relu_134;
assign relu_134[15:0] = (bias_add_134[31]==0) ? ((bias_add_134<3'd6) ? {{bias_add_134[31],bias_add_134[17:3]}} :'d6) : '0;
logic [15:0] relu_135;
assign relu_135[15:0] = (bias_add_135[31]==0) ? ((bias_add_135<3'd6) ? {{bias_add_135[31],bias_add_135[17:3]}} :'d6) : '0;
logic [15:0] relu_136;
assign relu_136[15:0] = (bias_add_136[31]==0) ? ((bias_add_136<3'd6) ? {{bias_add_136[31],bias_add_136[17:3]}} :'d6) : '0;
logic [15:0] relu_137;
assign relu_137[15:0] = (bias_add_137[31]==0) ? ((bias_add_137<3'd6) ? {{bias_add_137[31],bias_add_137[17:3]}} :'d6) : '0;
logic [15:0] relu_138;
assign relu_138[15:0] = (bias_add_138[31]==0) ? ((bias_add_138<3'd6) ? {{bias_add_138[31],bias_add_138[17:3]}} :'d6) : '0;
logic [15:0] relu_139;
assign relu_139[15:0] = (bias_add_139[31]==0) ? ((bias_add_139<3'd6) ? {{bias_add_139[31],bias_add_139[17:3]}} :'d6) : '0;
logic [15:0] relu_140;
assign relu_140[15:0] = (bias_add_140[31]==0) ? ((bias_add_140<3'd6) ? {{bias_add_140[31],bias_add_140[17:3]}} :'d6) : '0;
logic [15:0] relu_141;
assign relu_141[15:0] = (bias_add_141[31]==0) ? ((bias_add_141<3'd6) ? {{bias_add_141[31],bias_add_141[17:3]}} :'d6) : '0;
logic [15:0] relu_142;
assign relu_142[15:0] = (bias_add_142[31]==0) ? ((bias_add_142<3'd6) ? {{bias_add_142[31],bias_add_142[17:3]}} :'d6) : '0;
logic [15:0] relu_143;
assign relu_143[15:0] = (bias_add_143[31]==0) ? ((bias_add_143<3'd6) ? {{bias_add_143[31],bias_add_143[17:3]}} :'d6) : '0;
logic [15:0] relu_144;
assign relu_144[15:0] = (bias_add_144[31]==0) ? ((bias_add_144<3'd6) ? {{bias_add_144[31],bias_add_144[17:3]}} :'d6) : '0;
logic [15:0] relu_145;
assign relu_145[15:0] = (bias_add_145[31]==0) ? ((bias_add_145<3'd6) ? {{bias_add_145[31],bias_add_145[17:3]}} :'d6) : '0;
logic [15:0] relu_146;
assign relu_146[15:0] = (bias_add_146[31]==0) ? ((bias_add_146<3'd6) ? {{bias_add_146[31],bias_add_146[17:3]}} :'d6) : '0;
logic [15:0] relu_147;
assign relu_147[15:0] = (bias_add_147[31]==0) ? ((bias_add_147<3'd6) ? {{bias_add_147[31],bias_add_147[17:3]}} :'d6) : '0;
logic [15:0] relu_148;
assign relu_148[15:0] = (bias_add_148[31]==0) ? ((bias_add_148<3'd6) ? {{bias_add_148[31],bias_add_148[17:3]}} :'d6) : '0;
logic [15:0] relu_149;
assign relu_149[15:0] = (bias_add_149[31]==0) ? ((bias_add_149<3'd6) ? {{bias_add_149[31],bias_add_149[17:3]}} :'d6) : '0;
logic [15:0] relu_150;
assign relu_150[15:0] = (bias_add_150[31]==0) ? ((bias_add_150<3'd6) ? {{bias_add_150[31],bias_add_150[17:3]}} :'d6) : '0;
logic [15:0] relu_151;
assign relu_151[15:0] = (bias_add_151[31]==0) ? ((bias_add_151<3'd6) ? {{bias_add_151[31],bias_add_151[17:3]}} :'d6) : '0;
logic [15:0] relu_152;
assign relu_152[15:0] = (bias_add_152[31]==0) ? ((bias_add_152<3'd6) ? {{bias_add_152[31],bias_add_152[17:3]}} :'d6) : '0;
logic [15:0] relu_153;
assign relu_153[15:0] = (bias_add_153[31]==0) ? ((bias_add_153<3'd6) ? {{bias_add_153[31],bias_add_153[17:3]}} :'d6) : '0;
logic [15:0] relu_154;
assign relu_154[15:0] = (bias_add_154[31]==0) ? ((bias_add_154<3'd6) ? {{bias_add_154[31],bias_add_154[17:3]}} :'d6) : '0;
logic [15:0] relu_155;
assign relu_155[15:0] = (bias_add_155[31]==0) ? ((bias_add_155<3'd6) ? {{bias_add_155[31],bias_add_155[17:3]}} :'d6) : '0;
logic [15:0] relu_156;
assign relu_156[15:0] = (bias_add_156[31]==0) ? ((bias_add_156<3'd6) ? {{bias_add_156[31],bias_add_156[17:3]}} :'d6) : '0;
logic [15:0] relu_157;
assign relu_157[15:0] = (bias_add_157[31]==0) ? ((bias_add_157<3'd6) ? {{bias_add_157[31],bias_add_157[17:3]}} :'d6) : '0;
logic [15:0] relu_158;
assign relu_158[15:0] = (bias_add_158[31]==0) ? ((bias_add_158<3'd6) ? {{bias_add_158[31],bias_add_158[17:3]}} :'d6) : '0;
logic [15:0] relu_159;
assign relu_159[15:0] = (bias_add_159[31]==0) ? ((bias_add_159<3'd6) ? {{bias_add_159[31],bias_add_159[17:3]}} :'d6) : '0;
logic [15:0] relu_160;
assign relu_160[15:0] = (bias_add_160[31]==0) ? ((bias_add_160<3'd6) ? {{bias_add_160[31],bias_add_160[17:3]}} :'d6) : '0;
logic [15:0] relu_161;
assign relu_161[15:0] = (bias_add_161[31]==0) ? ((bias_add_161<3'd6) ? {{bias_add_161[31],bias_add_161[17:3]}} :'d6) : '0;
logic [15:0] relu_162;
assign relu_162[15:0] = (bias_add_162[31]==0) ? ((bias_add_162<3'd6) ? {{bias_add_162[31],bias_add_162[17:3]}} :'d6) : '0;
logic [15:0] relu_163;
assign relu_163[15:0] = (bias_add_163[31]==0) ? ((bias_add_163<3'd6) ? {{bias_add_163[31],bias_add_163[17:3]}} :'d6) : '0;
logic [15:0] relu_164;
assign relu_164[15:0] = (bias_add_164[31]==0) ? ((bias_add_164<3'd6) ? {{bias_add_164[31],bias_add_164[17:3]}} :'d6) : '0;
logic [15:0] relu_165;
assign relu_165[15:0] = (bias_add_165[31]==0) ? ((bias_add_165<3'd6) ? {{bias_add_165[31],bias_add_165[17:3]}} :'d6) : '0;
logic [15:0] relu_166;
assign relu_166[15:0] = (bias_add_166[31]==0) ? ((bias_add_166<3'd6) ? {{bias_add_166[31],bias_add_166[17:3]}} :'d6) : '0;
logic [15:0] relu_167;
assign relu_167[15:0] = (bias_add_167[31]==0) ? ((bias_add_167<3'd6) ? {{bias_add_167[31],bias_add_167[17:3]}} :'d6) : '0;
logic [15:0] relu_168;
assign relu_168[15:0] = (bias_add_168[31]==0) ? ((bias_add_168<3'd6) ? {{bias_add_168[31],bias_add_168[17:3]}} :'d6) : '0;
logic [15:0] relu_169;
assign relu_169[15:0] = (bias_add_169[31]==0) ? ((bias_add_169<3'd6) ? {{bias_add_169[31],bias_add_169[17:3]}} :'d6) : '0;
logic [15:0] relu_170;
assign relu_170[15:0] = (bias_add_170[31]==0) ? ((bias_add_170<3'd6) ? {{bias_add_170[31],bias_add_170[17:3]}} :'d6) : '0;
logic [15:0] relu_171;
assign relu_171[15:0] = (bias_add_171[31]==0) ? ((bias_add_171<3'd6) ? {{bias_add_171[31],bias_add_171[17:3]}} :'d6) : '0;
logic [15:0] relu_172;
assign relu_172[15:0] = (bias_add_172[31]==0) ? ((bias_add_172<3'd6) ? {{bias_add_172[31],bias_add_172[17:3]}} :'d6) : '0;
logic [15:0] relu_173;
assign relu_173[15:0] = (bias_add_173[31]==0) ? ((bias_add_173<3'd6) ? {{bias_add_173[31],bias_add_173[17:3]}} :'d6) : '0;
logic [15:0] relu_174;
assign relu_174[15:0] = (bias_add_174[31]==0) ? ((bias_add_174<3'd6) ? {{bias_add_174[31],bias_add_174[17:3]}} :'d6) : '0;
logic [15:0] relu_175;
assign relu_175[15:0] = (bias_add_175[31]==0) ? ((bias_add_175<3'd6) ? {{bias_add_175[31],bias_add_175[17:3]}} :'d6) : '0;
logic [15:0] relu_176;
assign relu_176[15:0] = (bias_add_176[31]==0) ? ((bias_add_176<3'd6) ? {{bias_add_176[31],bias_add_176[17:3]}} :'d6) : '0;
logic [15:0] relu_177;
assign relu_177[15:0] = (bias_add_177[31]==0) ? ((bias_add_177<3'd6) ? {{bias_add_177[31],bias_add_177[17:3]}} :'d6) : '0;
logic [15:0] relu_178;
assign relu_178[15:0] = (bias_add_178[31]==0) ? ((bias_add_178<3'd6) ? {{bias_add_178[31],bias_add_178[17:3]}} :'d6) : '0;
logic [15:0] relu_179;
assign relu_179[15:0] = (bias_add_179[31]==0) ? ((bias_add_179<3'd6) ? {{bias_add_179[31],bias_add_179[17:3]}} :'d6) : '0;
logic [15:0] relu_180;
assign relu_180[15:0] = (bias_add_180[31]==0) ? ((bias_add_180<3'd6) ? {{bias_add_180[31],bias_add_180[17:3]}} :'d6) : '0;
logic [15:0] relu_181;
assign relu_181[15:0] = (bias_add_181[31]==0) ? ((bias_add_181<3'd6) ? {{bias_add_181[31],bias_add_181[17:3]}} :'d6) : '0;
logic [15:0] relu_182;
assign relu_182[15:0] = (bias_add_182[31]==0) ? ((bias_add_182<3'd6) ? {{bias_add_182[31],bias_add_182[17:3]}} :'d6) : '0;
logic [15:0] relu_183;
assign relu_183[15:0] = (bias_add_183[31]==0) ? ((bias_add_183<3'd6) ? {{bias_add_183[31],bias_add_183[17:3]}} :'d6) : '0;
logic [15:0] relu_184;
assign relu_184[15:0] = (bias_add_184[31]==0) ? ((bias_add_184<3'd6) ? {{bias_add_184[31],bias_add_184[17:3]}} :'d6) : '0;
logic [15:0] relu_185;
assign relu_185[15:0] = (bias_add_185[31]==0) ? ((bias_add_185<3'd6) ? {{bias_add_185[31],bias_add_185[17:3]}} :'d6) : '0;
logic [15:0] relu_186;
assign relu_186[15:0] = (bias_add_186[31]==0) ? ((bias_add_186<3'd6) ? {{bias_add_186[31],bias_add_186[17:3]}} :'d6) : '0;
logic [15:0] relu_187;
assign relu_187[15:0] = (bias_add_187[31]==0) ? ((bias_add_187<3'd6) ? {{bias_add_187[31],bias_add_187[17:3]}} :'d6) : '0;
logic [15:0] relu_188;
assign relu_188[15:0] = (bias_add_188[31]==0) ? ((bias_add_188<3'd6) ? {{bias_add_188[31],bias_add_188[17:3]}} :'d6) : '0;
logic [15:0] relu_189;
assign relu_189[15:0] = (bias_add_189[31]==0) ? ((bias_add_189<3'd6) ? {{bias_add_189[31],bias_add_189[17:3]}} :'d6) : '0;
logic [15:0] relu_190;
assign relu_190[15:0] = (bias_add_190[31]==0) ? ((bias_add_190<3'd6) ? {{bias_add_190[31],bias_add_190[17:3]}} :'d6) : '0;
logic [15:0] relu_191;
assign relu_191[15:0] = (bias_add_191[31]==0) ? ((bias_add_191<3'd6) ? {{bias_add_191[31],bias_add_191[17:3]}} :'d6) : '0;
logic [15:0] relu_192;
assign relu_192[15:0] = (bias_add_192[31]==0) ? ((bias_add_192<3'd6) ? {{bias_add_192[31],bias_add_192[17:3]}} :'d6) : '0;
logic [15:0] relu_193;
assign relu_193[15:0] = (bias_add_193[31]==0) ? ((bias_add_193<3'd6) ? {{bias_add_193[31],bias_add_193[17:3]}} :'d6) : '0;
logic [15:0] relu_194;
assign relu_194[15:0] = (bias_add_194[31]==0) ? ((bias_add_194<3'd6) ? {{bias_add_194[31],bias_add_194[17:3]}} :'d6) : '0;
logic [15:0] relu_195;
assign relu_195[15:0] = (bias_add_195[31]==0) ? ((bias_add_195<3'd6) ? {{bias_add_195[31],bias_add_195[17:3]}} :'d6) : '0;
logic [15:0] relu_196;
assign relu_196[15:0] = (bias_add_196[31]==0) ? ((bias_add_196<3'd6) ? {{bias_add_196[31],bias_add_196[17:3]}} :'d6) : '0;
logic [15:0] relu_197;
assign relu_197[15:0] = (bias_add_197[31]==0) ? ((bias_add_197<3'd6) ? {{bias_add_197[31],bias_add_197[17:3]}} :'d6) : '0;
logic [15:0] relu_198;
assign relu_198[15:0] = (bias_add_198[31]==0) ? ((bias_add_198<3'd6) ? {{bias_add_198[31],bias_add_198[17:3]}} :'d6) : '0;
logic [15:0] relu_199;
assign relu_199[15:0] = (bias_add_199[31]==0) ? ((bias_add_199<3'd6) ? {{bias_add_199[31],bias_add_199[17:3]}} :'d6) : '0;
logic [15:0] relu_200;
assign relu_200[15:0] = (bias_add_200[31]==0) ? ((bias_add_200<3'd6) ? {{bias_add_200[31],bias_add_200[17:3]}} :'d6) : '0;
logic [15:0] relu_201;
assign relu_201[15:0] = (bias_add_201[31]==0) ? ((bias_add_201<3'd6) ? {{bias_add_201[31],bias_add_201[17:3]}} :'d6) : '0;
logic [15:0] relu_202;
assign relu_202[15:0] = (bias_add_202[31]==0) ? ((bias_add_202<3'd6) ? {{bias_add_202[31],bias_add_202[17:3]}} :'d6) : '0;
logic [15:0] relu_203;
assign relu_203[15:0] = (bias_add_203[31]==0) ? ((bias_add_203<3'd6) ? {{bias_add_203[31],bias_add_203[17:3]}} :'d6) : '0;
logic [15:0] relu_204;
assign relu_204[15:0] = (bias_add_204[31]==0) ? ((bias_add_204<3'd6) ? {{bias_add_204[31],bias_add_204[17:3]}} :'d6) : '0;
logic [15:0] relu_205;
assign relu_205[15:0] = (bias_add_205[31]==0) ? ((bias_add_205<3'd6) ? {{bias_add_205[31],bias_add_205[17:3]}} :'d6) : '0;
logic [15:0] relu_206;
assign relu_206[15:0] = (bias_add_206[31]==0) ? ((bias_add_206<3'd6) ? {{bias_add_206[31],bias_add_206[17:3]}} :'d6) : '0;
logic [15:0] relu_207;
assign relu_207[15:0] = (bias_add_207[31]==0) ? ((bias_add_207<3'd6) ? {{bias_add_207[31],bias_add_207[17:3]}} :'d6) : '0;
logic [15:0] relu_208;
assign relu_208[15:0] = (bias_add_208[31]==0) ? ((bias_add_208<3'd6) ? {{bias_add_208[31],bias_add_208[17:3]}} :'d6) : '0;
logic [15:0] relu_209;
assign relu_209[15:0] = (bias_add_209[31]==0) ? ((bias_add_209<3'd6) ? {{bias_add_209[31],bias_add_209[17:3]}} :'d6) : '0;
logic [15:0] relu_210;
assign relu_210[15:0] = (bias_add_210[31]==0) ? ((bias_add_210<3'd6) ? {{bias_add_210[31],bias_add_210[17:3]}} :'d6) : '0;
logic [15:0] relu_211;
assign relu_211[15:0] = (bias_add_211[31]==0) ? ((bias_add_211<3'd6) ? {{bias_add_211[31],bias_add_211[17:3]}} :'d6) : '0;
logic [15:0] relu_212;
assign relu_212[15:0] = (bias_add_212[31]==0) ? ((bias_add_212<3'd6) ? {{bias_add_212[31],bias_add_212[17:3]}} :'d6) : '0;
logic [15:0] relu_213;
assign relu_213[15:0] = (bias_add_213[31]==0) ? ((bias_add_213<3'd6) ? {{bias_add_213[31],bias_add_213[17:3]}} :'d6) : '0;
logic [15:0] relu_214;
assign relu_214[15:0] = (bias_add_214[31]==0) ? ((bias_add_214<3'd6) ? {{bias_add_214[31],bias_add_214[17:3]}} :'d6) : '0;
logic [15:0] relu_215;
assign relu_215[15:0] = (bias_add_215[31]==0) ? ((bias_add_215<3'd6) ? {{bias_add_215[31],bias_add_215[17:3]}} :'d6) : '0;
logic [15:0] relu_216;
assign relu_216[15:0] = (bias_add_216[31]==0) ? ((bias_add_216<3'd6) ? {{bias_add_216[31],bias_add_216[17:3]}} :'d6) : '0;
logic [15:0] relu_217;
assign relu_217[15:0] = (bias_add_217[31]==0) ? ((bias_add_217<3'd6) ? {{bias_add_217[31],bias_add_217[17:3]}} :'d6) : '0;
logic [15:0] relu_218;
assign relu_218[15:0] = (bias_add_218[31]==0) ? ((bias_add_218<3'd6) ? {{bias_add_218[31],bias_add_218[17:3]}} :'d6) : '0;
logic [15:0] relu_219;
assign relu_219[15:0] = (bias_add_219[31]==0) ? ((bias_add_219<3'd6) ? {{bias_add_219[31],bias_add_219[17:3]}} :'d6) : '0;
logic [15:0] relu_220;
assign relu_220[15:0] = (bias_add_220[31]==0) ? ((bias_add_220<3'd6) ? {{bias_add_220[31],bias_add_220[17:3]}} :'d6) : '0;
logic [15:0] relu_221;
assign relu_221[15:0] = (bias_add_221[31]==0) ? ((bias_add_221<3'd6) ? {{bias_add_221[31],bias_add_221[17:3]}} :'d6) : '0;
logic [15:0] relu_222;
assign relu_222[15:0] = (bias_add_222[31]==0) ? ((bias_add_222<3'd6) ? {{bias_add_222[31],bias_add_222[17:3]}} :'d6) : '0;
logic [15:0] relu_223;
assign relu_223[15:0] = (bias_add_223[31]==0) ? ((bias_add_223<3'd6) ? {{bias_add_223[31],bias_add_223[17:3]}} :'d6) : '0;
logic [15:0] relu_224;
assign relu_224[15:0] = (bias_add_224[31]==0) ? ((bias_add_224<3'd6) ? {{bias_add_224[31],bias_add_224[17:3]}} :'d6) : '0;
logic [15:0] relu_225;
assign relu_225[15:0] = (bias_add_225[31]==0) ? ((bias_add_225<3'd6) ? {{bias_add_225[31],bias_add_225[17:3]}} :'d6) : '0;
logic [15:0] relu_226;
assign relu_226[15:0] = (bias_add_226[31]==0) ? ((bias_add_226<3'd6) ? {{bias_add_226[31],bias_add_226[17:3]}} :'d6) : '0;
logic [15:0] relu_227;
assign relu_227[15:0] = (bias_add_227[31]==0) ? ((bias_add_227<3'd6) ? {{bias_add_227[31],bias_add_227[17:3]}} :'d6) : '0;
logic [15:0] relu_228;
assign relu_228[15:0] = (bias_add_228[31]==0) ? ((bias_add_228<3'd6) ? {{bias_add_228[31],bias_add_228[17:3]}} :'d6) : '0;
logic [15:0] relu_229;
assign relu_229[15:0] = (bias_add_229[31]==0) ? ((bias_add_229<3'd6) ? {{bias_add_229[31],bias_add_229[17:3]}} :'d6) : '0;
logic [15:0] relu_230;
assign relu_230[15:0] = (bias_add_230[31]==0) ? ((bias_add_230<3'd6) ? {{bias_add_230[31],bias_add_230[17:3]}} :'d6) : '0;
logic [15:0] relu_231;
assign relu_231[15:0] = (bias_add_231[31]==0) ? ((bias_add_231<3'd6) ? {{bias_add_231[31],bias_add_231[17:3]}} :'d6) : '0;
logic [15:0] relu_232;
assign relu_232[15:0] = (bias_add_232[31]==0) ? ((bias_add_232<3'd6) ? {{bias_add_232[31],bias_add_232[17:3]}} :'d6) : '0;
logic [15:0] relu_233;
assign relu_233[15:0] = (bias_add_233[31]==0) ? ((bias_add_233<3'd6) ? {{bias_add_233[31],bias_add_233[17:3]}} :'d6) : '0;
logic [15:0] relu_234;
assign relu_234[15:0] = (bias_add_234[31]==0) ? ((bias_add_234<3'd6) ? {{bias_add_234[31],bias_add_234[17:3]}} :'d6) : '0;
logic [15:0] relu_235;
assign relu_235[15:0] = (bias_add_235[31]==0) ? ((bias_add_235<3'd6) ? {{bias_add_235[31],bias_add_235[17:3]}} :'d6) : '0;
logic [15:0] relu_236;
assign relu_236[15:0] = (bias_add_236[31]==0) ? ((bias_add_236<3'd6) ? {{bias_add_236[31],bias_add_236[17:3]}} :'d6) : '0;
logic [15:0] relu_237;
assign relu_237[15:0] = (bias_add_237[31]==0) ? ((bias_add_237<3'd6) ? {{bias_add_237[31],bias_add_237[17:3]}} :'d6) : '0;
logic [15:0] relu_238;
assign relu_238[15:0] = (bias_add_238[31]==0) ? ((bias_add_238<3'd6) ? {{bias_add_238[31],bias_add_238[17:3]}} :'d6) : '0;
logic [15:0] relu_239;
assign relu_239[15:0] = (bias_add_239[31]==0) ? ((bias_add_239<3'd6) ? {{bias_add_239[31],bias_add_239[17:3]}} :'d6) : '0;
logic [15:0] relu_240;
assign relu_240[15:0] = (bias_add_240[31]==0) ? ((bias_add_240<3'd6) ? {{bias_add_240[31],bias_add_240[17:3]}} :'d6) : '0;
logic [15:0] relu_241;
assign relu_241[15:0] = (bias_add_241[31]==0) ? ((bias_add_241<3'd6) ? {{bias_add_241[31],bias_add_241[17:3]}} :'d6) : '0;
logic [15:0] relu_242;
assign relu_242[15:0] = (bias_add_242[31]==0) ? ((bias_add_242<3'd6) ? {{bias_add_242[31],bias_add_242[17:3]}} :'d6) : '0;
logic [15:0] relu_243;
assign relu_243[15:0] = (bias_add_243[31]==0) ? ((bias_add_243<3'd6) ? {{bias_add_243[31],bias_add_243[17:3]}} :'d6) : '0;
logic [15:0] relu_244;
assign relu_244[15:0] = (bias_add_244[31]==0) ? ((bias_add_244<3'd6) ? {{bias_add_244[31],bias_add_244[17:3]}} :'d6) : '0;
logic [15:0] relu_245;
assign relu_245[15:0] = (bias_add_245[31]==0) ? ((bias_add_245<3'd6) ? {{bias_add_245[31],bias_add_245[17:3]}} :'d6) : '0;
logic [15:0] relu_246;
assign relu_246[15:0] = (bias_add_246[31]==0) ? ((bias_add_246<3'd6) ? {{bias_add_246[31],bias_add_246[17:3]}} :'d6) : '0;
logic [15:0] relu_247;
assign relu_247[15:0] = (bias_add_247[31]==0) ? ((bias_add_247<3'd6) ? {{bias_add_247[31],bias_add_247[17:3]}} :'d6) : '0;
logic [15:0] relu_248;
assign relu_248[15:0] = (bias_add_248[31]==0) ? ((bias_add_248<3'd6) ? {{bias_add_248[31],bias_add_248[17:3]}} :'d6) : '0;
logic [15:0] relu_249;
assign relu_249[15:0] = (bias_add_249[31]==0) ? ((bias_add_249<3'd6) ? {{bias_add_249[31],bias_add_249[17:3]}} :'d6) : '0;
logic [15:0] relu_250;
assign relu_250[15:0] = (bias_add_250[31]==0) ? ((bias_add_250<3'd6) ? {{bias_add_250[31],bias_add_250[17:3]}} :'d6) : '0;
logic [15:0] relu_251;
assign relu_251[15:0] = (bias_add_251[31]==0) ? ((bias_add_251<3'd6) ? {{bias_add_251[31],bias_add_251[17:3]}} :'d6) : '0;
logic [15:0] relu_252;
assign relu_252[15:0] = (bias_add_252[31]==0) ? ((bias_add_252<3'd6) ? {{bias_add_252[31],bias_add_252[17:3]}} :'d6) : '0;
logic [15:0] relu_253;
assign relu_253[15:0] = (bias_add_253[31]==0) ? ((bias_add_253<3'd6) ? {{bias_add_253[31],bias_add_253[17:3]}} :'d6) : '0;
logic [15:0] relu_254;
assign relu_254[15:0] = (bias_add_254[31]==0) ? ((bias_add_254<3'd6) ? {{bias_add_254[31],bias_add_254[17:3]}} :'d6) : '0;
logic [15:0] relu_255;
assign relu_255[15:0] = (bias_add_255[31]==0) ? ((bias_add_255<3'd6) ? {{bias_add_255[31],bias_add_255[17:3]}} :'d6) : '0;

assign output_act = {
	relu_255,
	relu_254,
	relu_253,
	relu_252,
	relu_251,
	relu_250,
	relu_249,
	relu_248,
	relu_247,
	relu_246,
	relu_245,
	relu_244,
	relu_243,
	relu_242,
	relu_241,
	relu_240,
	relu_239,
	relu_238,
	relu_237,
	relu_236,
	relu_235,
	relu_234,
	relu_233,
	relu_232,
	relu_231,
	relu_230,
	relu_229,
	relu_228,
	relu_227,
	relu_226,
	relu_225,
	relu_224,
	relu_223,
	relu_222,
	relu_221,
	relu_220,
	relu_219,
	relu_218,
	relu_217,
	relu_216,
	relu_215,
	relu_214,
	relu_213,
	relu_212,
	relu_211,
	relu_210,
	relu_209,
	relu_208,
	relu_207,
	relu_206,
	relu_205,
	relu_204,
	relu_203,
	relu_202,
	relu_201,
	relu_200,
	relu_199,
	relu_198,
	relu_197,
	relu_196,
	relu_195,
	relu_194,
	relu_193,
	relu_192,
	relu_191,
	relu_190,
	relu_189,
	relu_188,
	relu_187,
	relu_186,
	relu_185,
	relu_184,
	relu_183,
	relu_182,
	relu_181,
	relu_180,
	relu_179,
	relu_178,
	relu_177,
	relu_176,
	relu_175,
	relu_174,
	relu_173,
	relu_172,
	relu_171,
	relu_170,
	relu_169,
	relu_168,
	relu_167,
	relu_166,
	relu_165,
	relu_164,
	relu_163,
	relu_162,
	relu_161,
	relu_160,
	relu_159,
	relu_158,
	relu_157,
	relu_156,
	relu_155,
	relu_154,
	relu_153,
	relu_152,
	relu_151,
	relu_150,
	relu_149,
	relu_148,
	relu_147,
	relu_146,
	relu_145,
	relu_144,
	relu_143,
	relu_142,
	relu_141,
	relu_140,
	relu_139,
	relu_138,
	relu_137,
	relu_136,
	relu_135,
	relu_134,
	relu_133,
	relu_132,
	relu_131,
	relu_130,
	relu_129,
	relu_128,
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
